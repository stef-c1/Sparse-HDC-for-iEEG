module dense_skel # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125, //0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer LBP_LENGTH = 6,
    parameter integer NB_CLASSES = 2,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk_i,
    input  arst_n_in,
    input  [LBP_LENGTH-1:0] LBP_codes63,
    input  [LBP_LENGTH-1:0] LBP_codes62,
    input  [LBP_LENGTH-1:0] LBP_codes61,
    input  [LBP_LENGTH-1:0] LBP_codes60,
    input  [LBP_LENGTH-1:0] LBP_codes59,
    input  [LBP_LENGTH-1:0] LBP_codes58,
    input  [LBP_LENGTH-1:0] LBP_codes57,
    input  [LBP_LENGTH-1:0] LBP_codes56,
    input  [LBP_LENGTH-1:0] LBP_codes55,
    input  [LBP_LENGTH-1:0] LBP_codes54,
    input  [LBP_LENGTH-1:0] LBP_codes53,
    input  [LBP_LENGTH-1:0] LBP_codes52,
    input  [LBP_LENGTH-1:0] LBP_codes51,
    input  [LBP_LENGTH-1:0] LBP_codes50,
    input  [LBP_LENGTH-1:0] LBP_codes49,
    input  [LBP_LENGTH-1:0] LBP_codes48,
    input  [LBP_LENGTH-1:0] LBP_codes47,
    input  [LBP_LENGTH-1:0] LBP_codes46,
    input  [LBP_LENGTH-1:0] LBP_codes45,
    input  [LBP_LENGTH-1:0] LBP_codes44,
    input  [LBP_LENGTH-1:0] LBP_codes43,
    input  [LBP_LENGTH-1:0] LBP_codes42,
    input  [LBP_LENGTH-1:0] LBP_codes41,
    input  [LBP_LENGTH-1:0] LBP_codes40,
    input  [LBP_LENGTH-1:0] LBP_codes39,
    input  [LBP_LENGTH-1:0] LBP_codes38,
    input  [LBP_LENGTH-1:0] LBP_codes37,
    input  [LBP_LENGTH-1:0] LBP_codes36,
    input  [LBP_LENGTH-1:0] LBP_codes35,
    input  [LBP_LENGTH-1:0] LBP_codes34,
    input  [LBP_LENGTH-1:0] LBP_codes33,
    input  [LBP_LENGTH-1:0] LBP_codes32,
    input  [LBP_LENGTH-1:0] LBP_codes31,
    input  [LBP_LENGTH-1:0] LBP_codes30,
    input  [LBP_LENGTH-1:0] LBP_codes29,
    input  [LBP_LENGTH-1:0] LBP_codes28,
    input  [LBP_LENGTH-1:0] LBP_codes27,
    input  [LBP_LENGTH-1:0] LBP_codes26,
    input  [LBP_LENGTH-1:0] LBP_codes25,
    input  [LBP_LENGTH-1:0] LBP_codes24,
    input  [LBP_LENGTH-1:0] LBP_codes23,
    input  [LBP_LENGTH-1:0] LBP_codes22,
    input  [LBP_LENGTH-1:0] LBP_codes21,
    input  [LBP_LENGTH-1:0] LBP_codes20,
    input  [LBP_LENGTH-1:0] LBP_codes19,
    input  [LBP_LENGTH-1:0] LBP_codes18,
    input  [LBP_LENGTH-1:0] LBP_codes17,
    input  [LBP_LENGTH-1:0] LBP_codes16,
    input  [LBP_LENGTH-1:0] LBP_codes15,
    input  [LBP_LENGTH-1:0] LBP_codes14,
    input  [LBP_LENGTH-1:0] LBP_codes13,
    input  [LBP_LENGTH-1:0] LBP_codes12,
    input  [LBP_LENGTH-1:0] LBP_codes11,
    input  [LBP_LENGTH-1:0] LBP_codes10,
    input  [LBP_LENGTH-1:0] LBP_codes9,
    input  [LBP_LENGTH-1:0] LBP_codes8,
    input  [LBP_LENGTH-1:0] LBP_codes7,
    input  [LBP_LENGTH-1:0] LBP_codes6,
    input  [LBP_LENGTH-1:0] LBP_codes5,
    input  [LBP_LENGTH-1:0] LBP_codes4,
    input  [LBP_LENGTH-1:0] LBP_codes3,
    input  [LBP_LENGTH-1:0] LBP_codes2,
    input  [LBP_LENGTH-1:0] LBP_codes1,
    input  [LBP_LENGTH-1:0] LBP_codes0,
    input  [0:D-1] ictal_hv_in,
    input  [0:D-1] interictal_hv_in,
    output classification_ready,
    output [$clog2(NB_CLASSES)-1:0] classification,
    output send_next_LBP,
    output [$clog2(D):0] ictal_sim,
    output [$clog2(D):0] interictal_sim
);

//LBP_codes
logic [LBP_LENGTH-1:0] LBP_codes [E-1:0];
assign LBP_codes[63] = LBP_codes63;
assign LBP_codes[62] = LBP_codes62;
assign LBP_codes[61] = LBP_codes61;
assign LBP_codes[60] = LBP_codes60;
assign LBP_codes[59] = LBP_codes59;
assign LBP_codes[58] = LBP_codes58;
assign LBP_codes[57] = LBP_codes57;
assign LBP_codes[56] = LBP_codes56;
assign LBP_codes[55] = LBP_codes55;
assign LBP_codes[54] = LBP_codes54;
assign LBP_codes[53] = LBP_codes53;
assign LBP_codes[52] = LBP_codes52;
assign LBP_codes[51] = LBP_codes51;
assign LBP_codes[50] = LBP_codes50;
assign LBP_codes[49] = LBP_codes49;
assign LBP_codes[48] = LBP_codes48;
assign LBP_codes[47] = LBP_codes47;
assign LBP_codes[46] = LBP_codes46;
assign LBP_codes[45] = LBP_codes45;
assign LBP_codes[44] = LBP_codes44;
assign LBP_codes[43] = LBP_codes43;
assign LBP_codes[42] = LBP_codes42;
assign LBP_codes[41] = LBP_codes41;
assign LBP_codes[40] = LBP_codes40;
assign LBP_codes[39] = LBP_codes39;
assign LBP_codes[38] = LBP_codes38;
assign LBP_codes[37] = LBP_codes37;
assign LBP_codes[36] = LBP_codes36;
assign LBP_codes[35] = LBP_codes35;
assign LBP_codes[34] = LBP_codes34;
assign LBP_codes[33] = LBP_codes33;
assign LBP_codes[32] = LBP_codes32;
assign LBP_codes[31] = LBP_codes31;
assign LBP_codes[30] = LBP_codes30;
assign LBP_codes[29] = LBP_codes29;
assign LBP_codes[28] = LBP_codes28;
assign LBP_codes[27] = LBP_codes27;
assign LBP_codes[26] = LBP_codes26;
assign LBP_codes[25] = LBP_codes25;
assign LBP_codes[24] = LBP_codes24;
assign LBP_codes[23] = LBP_codes23;
assign LBP_codes[22] = LBP_codes22;
assign LBP_codes[21] = LBP_codes21;
assign LBP_codes[20] = LBP_codes20;
assign LBP_codes[19] = LBP_codes19;
assign LBP_codes[18] = LBP_codes18;
assign LBP_codes[17] = LBP_codes17;
assign LBP_codes[16] = LBP_codes16;
assign LBP_codes[15] = LBP_codes15;
assign LBP_codes[14] = LBP_codes14;
assign LBP_codes[13] = LBP_codes13;
assign LBP_codes[12] = LBP_codes12;
assign LBP_codes[11] = LBP_codes11;
assign LBP_codes[10] = LBP_codes10;
assign LBP_codes[9] = LBP_codes9;
assign LBP_codes[8] = LBP_codes8;
assign LBP_codes[7] = LBP_codes7;
assign LBP_codes[6] = LBP_codes6;
assign LBP_codes[5] = LBP_codes5;
assign LBP_codes[4] = LBP_codes4;
assign LBP_codes[3] = LBP_codes3;
assign LBP_codes[2] = LBP_codes2;
assign LBP_codes[1] = LBP_codes1;
assign LBP_codes[0] = LBP_codes0;



//signal that need next LBP_codes
assign send_next_LBP = 1;



logic [E-1:0][D-1:0] LBP_hvs;


logic [E-1:0][0:D-1] bind_outputs;


logic bundled_hv [0:D-1];


logic [0:D-1] result_hv;
logic [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time;
logic signed [4:0] counter_array [0:D-1];

logic [0:D-1] ictal_hv;
logic [0:D-1] interictal_hv;


assign ictal_hv = (arst_n_in) ? ictal_hv : ictal_hv_in;
assign interictal_hv = (arst_n_in) ? interictal_hv : interictal_hv_in;

//The Big Five
IM #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
IM_module (.clk_i(clk_i), .arst_n_in(arst_n_in), .LBP_codes(LBP_codes), .LBP_hvs(LBP_hvs));

BINDING #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BINDING_module (.LBP_hvs(LBP_hvs), .bind_outputs(bind_outputs));

BUNDLING_SPACE #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BUNDLING_SPACE_module (.clk_i(clk_i), .arst_n_in(arst_n_in), .bind_outputs(bind_outputs), .bundled_hv(bundled_hv));

BUNDLING_TIME #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .NB_TO_BUNDLE_IN_TIME(NB_TO_BUNDLE_IN_TIME), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BUNDLING_TIME_module (.clk_i(clk_i), .arst_n_in(arst_n_in), .bundled_hv(bundled_hv), .result_hv(result_hv), .counter_bund_time(counter_bund_time), .counter_array(counter_array));

SIMILARITY_SEARCH #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .NB_TO_BUNDLE_IN_TIME(NB_TO_BUNDLE_IN_TIME), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor), .NB_CLASSES(NB_CLASSES)) 
SIMILARITY_SEARCH_module (.clk_i(clk_i), .arst_n_in(arst_n_in), .result_hv(result_hv), .ictal_hv(ictal_hv), .interictal_hv(interictal_hv), .counter_bund_time(counter_bund_time), .classification(classification), .classification_ready(classification_ready), .ictal_sim(ictal_sim), .interictal_sim(interictal_sim));

endmodule


module IM # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk_i,
    input  arst_n_in,
    input  [LBP_LENGTH-1:0] LBP_codes [E-1:0],
    output logic [E-1:0][D-1:0] LBP_hvs
);

//IM
logic [2**(LBP_LENGTH)-1:0][D-1:0] IM;

assign IM[0] = 1024'b1000010011011001011100101011000011101001000110001011100001110110011100010111101001010100011101101010110111010011100000001011001001000010100101101110101000101001010110001100001111000111000010101110011010000100101001011101010110111101101101111001011011001111111010010101010100000011010011100111011010110111010101000000100100001011000001101111001010000010010101100110000011101001101101111010110001101111000010101100101010100010111100111010001001001101100010111000010100110000001010010010101111001110101100100101001110111101011111111000100011100000101101011101010010100100110101111111110010100010000111111011100001111010001111100010011110000101101000001100000000101110010011010111001110101011111101000000100101001100110101101010101010001000101001100100010101110110000111000110010011101101001011001111110011100000000101010001100111000110110001101110111011010001111101001100110111111000111000111111101000101011000000100100100001011101011011011110010010101000011110101111001000110111011011101011110010000100010000000110101011101111;
assign IM[1] = 1024'b1000110011001101110100111001111001000101000111011001110100001010100110100001000001101010001100001000010100111010001000000110001111000010010111100010010101010001101011010011110111010101100011001011100111000111101001101100011000011100111010011000100110000010011110101010111001010000101100100000100111000101000001000111100011110110100111100100011010110011010101010001000111000110100110100111111001010011101011101010010000111100110101000000000010110110001000101100110011111001100111001100011110011111110110100001100111110100000000001000111001101001110011010011101111100010001000011001001011010011000001110100001111011100101111000011000101011101110010110100011011000011001100010111100001111111000011100010101110001110101111110001100000110001010100100011000111001111101100001110111011111011100100001100111001011010100101001011011110011001000010011110000111111101001101111100010101101010101111110011101000011001011100101001000111000100011110010110111111111101110001100000110100011110011101111100111111110101100000010010010101011001;
assign IM[2] = 1024'b0000000101111011111000110110010110001101101110100010000101110000101110001111110111011110101011001010011100011101111001110001110000101010011001000111100001111010110111111111010100111110001000001000011011100010011110011101000001110101101011000011011000101001000111101100010010010111110101000100100101011011010100010001101100010000010011100000110101100011101001011110001111101000111100110010000010110100111001000101001010000010000101011010100010101010110100101100011001111111110000000111000101000010011000110011001101011111011000110011111110010011001001011011001101010101111001000011110111101010000010011010111101001111010000010001100000000100110010010000101001100010101101101001111110101101011001001011010111110101101100010110001011101010000011111001011101110101011100010001010100001011100010111101100000101001001011100100000111111100101100000100010010010010111110001111001110101111111101011010111000001011000100110111101100111111000101010111011100010110010000001001111100101000101000001000000101111001110110110110000011111101;
assign IM[3] = 1024'b1011011001011010100000010011001011011011100110111101011010011001010010110101010000001001111000000110101101101100001110100111111101101110111010100011001010010010001000001010110011010100100111000001101100001101001011010011110000100011011001000001010000110110000110111110100110001011110100100100110000111010011101101110001010011100000010011101111101010110111100110010010111001001001011101101100100111010001111010010011110101101010110011000000011100000111101010001111011010110010100010111011100101010100110000101110111101010011100111101011001110111001110011010000101110100110100010011001100001001001111110001010110111011110001001100011011011111001110000101101111000110101110001100111110001011101010110011000101100100100100100010111101101011011100000011111111111000111110000100111001100100011000010010000110110011000011010000010001111001100001011111100001111110001101010010100100000100001100111010101000001001100100101101010000010110100111001010101101001010000011101100101101111011001110001110001111101000001101010001110001001101;
assign IM[4] = 1024'b0001111000010011010011101001001001100111101111110100111111100011011001001001001000100101000011101100110010110011001110100001010111011010110001010110001110000010110111101000001101010101100011001001110101110110110110010001111110000001111101111011011101100011101011110000110010010000001011011100011000000111111110010110111000111011110101111010011111110101000000111011001010110001101101100010011111010000100101110111001001000010111000100100101011100001011010000110011001110001110100010010100100000110110110010011000000000000101001110110101100110101101001001001010001101111111101101110011010101011110100001010001001000010110110101011100011001101110100110100011000111001011110000111001001010101100000010111101001110000101110101001001000001010110000010111011100101001111000110011100110011111100110100111101100001101000000111000101010010100101010110010000000110110010000110001111111110101101011111000100000011101001000111101100001100000000100000010110110001101110111000111001011111011110101000000111101111010100001010111011111101100;
assign IM[5] = 1024'b0100011001111111010101000101101100110110001101010011100111111101001100000111111001010000010000011011101010100100100101111101011011000000101001100000010000111000111100011110101010110100110000001101001001101110101111001000011000111001100001100100111011111110010110000000111001011001110101101000111001001001110111100000111100000011111101100101001001111001011011001110111111110110101110011111101110000100011101001101010111111111110011010001100000011001010101110011001110000111011111001100110110011001101111100000101000100000010010100101001111000110011110000010000011000101011110111001010000001101000011000100001111000010000010100011001101100101011000110100101010001100010000101100011000011111101011111111011000101000000001010100011010011100100110101001000000001101100010110011000000111000010100001101110110011011000101000101111100001111000111011101000111010011010001110001111001111101010110000001101011110001010101010000110100011101101111110100101110001101011111000011100000100110001111100111001001111110011000011010111111011110;
assign IM[6] = 1024'b1011111101111001010010100101110111001101001101001110010111010111101000101010010111100110011111100110110000011000110101000000110111011001100010010101111001000100010101000011010011000111100100101001000101101101100001001100111000000011011100000110000001101001010011011101000010111111100011000001011011001001101111011010101000110111101000110011010100101001001000111010000101010010111100001100110000100100010011000100110111100111100111010110000100110111001010000011100101000100100110010101100101110011000011000111100000101101101011100001001100111111010110011001010000110010111001011100101111011101110100001110100000101000011010010111100100101110010011011100101000010110011100100110100011110101111010000110110101101000110111101010010111110000001111110001101010100010010111110011110000110100111010011100001101111100111111010110010100101010011000101011111111111110011001111110000100000001101101011011100100111000111011011010101110001011001000010000101110011000101110010101101111100100000001000010011011010001101101011010010010010010;
assign IM[7] = 1024'b0111010010000101001011101001100101000010000101011010100010111001100001001001110011011100000111110101100100011010010101101110010100100110001011110111111001100110100111101011110101101001111001001111011100101110110110001000111001111000011010000011100011010101110010110000011110100110001011111111011000101110011101110011111110001001011100100001111101111110110101001111010100010101010100101100101001101011100110001000101011000101110010001010011001001001001011001100111001100001111000111101001111101010100101110101001001100110110111000110011101101010000001010111011101111100110001010100001010001011011011011001111000010011010010111100011000001001111011001010111000010000001011000000010000101100001101110000110110101010111100011110101110001101101111100010000010000011001101010011110010101110000011100110011000101101011000110001001010101101001100010001100001000100110110110110001110101110110011000001100000000110110111101000111100001011110111010111001000100001100101100111100101100000111011001110101100000101010111000000100011110110;
assign IM[8] = 1024'b0001001100000000011100010001010010110101000100001101110100111100100011010010011011111111010110001001000101111011101001011011111110110110110100001111111001011111000111110001111010011100011011011111001000010011011000111111001011111101000001110000111100001000001001010010001100000101100000000000100001011111010001110000110000001100000010001000010010001001111110101011001110101011110011110101110110011110110100110100001100111010001100100001001011001101100001111001110001011011101010110001100110101110110100000011111101101001100000010101100000110100111100101011001111100110011001010101000010100111100011111110001000011000001101111111101011000110111101111001100111100000110011110101111101001011111010000101001011110111110111000100000001100001010101110111101111000001100100100010110110000000110000001101001111101010100010111111111100100010111000100000010001011001011100000001110100010111101110000000111100001111110000110001100000100011111010010001100011111101110011001111001100010010111111100111000100100010101010111001001101110011;
assign IM[9] = 1024'b1011110110010100001010100100111010011011000100011011110000010111001011011101100010001010000101111011000111100000011111111010001000001111010010000000110111100010011101110001101101010010011101011101100000111000111010101001000100000101101100110101100010010000110101001110010000001000111000010011010111101000010011101111011110110001111000010101110100010100010101101101011100010001011111100001001001010111111110101110100001101111100110011110011001101011100100111001101110011011011001011001000010111000010011111011111111111111010111101101011000010110100001110111000111001110110010000110110000100001100100101011011100100100101001000010010101111110101010000000010110011101101010100111001100100011110011000111111111001010100000001101101010011001000111110001011111000001010110111000000000110100000000011001010110000111111111100110110001011000110100100101010100001000010100100111001001111001110011001011001111111101010101011011000101011111100000010010110000101010000010000011000111110011100111011110100001101000100110110000001111110111;
assign IM[10] = 1024'b0001101000010010001101011101000111000100111000111001011011011101110011100101101001011100001001011100100110010001000011110100111011011101001011100001100001100011001101011100010001111111111100110101011101111011100000101010111111000111110011010010001110101010000001110110101010111100001111101111111010000010001011101010100110011110111001101101011110100101110000010111000010001001111011111001111101011010111001110011111110101010011010001100111010010011111010100000001110011100100011110111111011101111110111001111110000111000011010100001101101001101110010110111110001011100010011010011111010001100001000001000100010100000011001001101101100011110111100000101100011001101001010001111011011100100001100101101010011111000100001101000110111000001011011101100100100101011000011111110001011111110010000111100001001101101010100000001110000000110101101110011001111110110011000011110000010000000000110000010000110101110011000011011000101010001110001010000011000010010000010000110010001010100001101001111010000001010010011001001111000101011;
assign IM[11] = 1024'b0111101011111001000111101111100101011101000010000111100111011110101100010110001011011100100110000011101010001101001100101111001101100011100001100001000001010101111011101101010011101001101111110011001100000101010101111110111101011111110000101001110110000110111010001110001111010110010011011010001010001100100010011111010011010010111101000001011111100110000100101110000100010110001100111100110110111110110010011110010101011011110100101100111010011101000101000111011010001010101001110100010010100100000011110101011110000010111100110010110010011100111111101000101101100110101110001100100110010101110101100001011101001000010100100110111110110100100000001100100000010100111110001100100111100000011010011110001100110010001001111110001010001011001000001010011001000111010010100000110111001110010101101000111011001010010001000000001000110000000011001001100011000111001101101111100111011110011100011011001111110010100001110110001101110000110000000111111111101001000101010000100010101110011010111100000110111001001111011000000110001100;
assign IM[12] = 1024'b1001001111001101101010001100111111111001111001001110111010001101001110000000011100001110001001011110001001101111010001111001100000111101010011100110000001000001000110101000001010110110111100011110000110001010111101101101000100110100101110111111100000001000101001011001000111010010110000000111010001001100100010100010111001010010001001110001000000000111011111010101011000111100000000100010110111010001011011010111110100110110011010110110001010111101011011111100101110110001111111011110011100110101001011101001010000110000100001101000101111001100011000101110000001011111111100100010101011010110101001111000000011111000110011100101000000100011111100111111100010101100111001110101011100111101010011010001101011001110011111010001101011001110011001000000100010000100110101001100101010111100001000000001000111110011010111011110100101110010110110000000101011000100001100101011000111001000001110000011011000111010001100110101110100001011011111001100111001011100101001111111011111010010100011101000010111110000111010110111011000111001;
assign IM[13] = 1024'b1011100100100101101011000101111001010100011100101011010000011011010100000110100001100101011011100100101100001111000111001101110101111111111011110110001011000101100001111011000000001000111100001100111100010010111011101111000011100001010110011100011000011001010111111011001000100011101101010101010100100000011001011101010000110000110100010110010000110100010101110001100100101100100001110001000000111101101101001010111000111010001001110101110010101000011111010101111110111001111000001111110001000110010010110011110101011110011110100100001111100010110101101010101011101000111010011000010000000101001101001011001001001011000010100011000000101010010101011101011001000001110100000001001011110010000001110110011011100000111000111011000010000111101010100000010100110101110011000100101111111111111011100000010101110001101110000100111101101101111010100011111110110000110111101000001010110101110111000000101001001011111110001011101010000011101011110111011011110010111001110100100011010000110001110011110110000101100110101100011111010011;
assign IM[14] = 1024'b1101110101011011110111100110111101011101011101001001001010010001100100111111011001001000001010010011110110010101111011111110100101111011100101111011100111000110100111101010100111001000000001101001011100100100110111100011111100001010000011000110010111010110100100110010110111001100010011100001101111100110000100000010100001000010000111111001000010100111001111010000100010101100001100111100011011110010011011001000110111001110100011011000011001001101000011111010000101101100010100101000110101000101001001010000100101010011100100000001001111011000011011111000011011010011101101010000111010001101110110110111110101011001110110111010110110101000011001010000000111000110101010001110100101001111110100001110101010000011110000010110011111001011100000010001000100110110011101100101110101000100111011101000101100000100100001011101110110110110000101100101000001010010000011110111010110000010111000100010010111100010001111100001001110010100101011101111111010011110011100000011001110011110110111011100101001110110110111010011100010100010;
assign IM[15] = 1024'b0110011000111110001000111000101010000100111100111100110010001000111100111111011001111110001101011100101111000100100001010101001010000000110100101011101010110001101011011000101111100100100101011001101011111010110100010011011010010110110100001010010110111011110011001010110111011101011110011110011001011010111001101010101000111100011010011010010111101001000010100111001011111100101100001100001100000010111001110000100100100101110000011101011111100110101111111010010111011010101000000100111010111100100010000100011101101000000010111000110010110000000111111011001000101110000011011010011010001011011000101001111000010011110111011000111101010111011011111100011100011111110101000001110100001000000011110001110101001001000100001110001101110111101011000011001000101111100100001110111011111101100000100111001100000011100010111110101110110110101101000100011110111100110001001100100000101001111111101101000000111001010001110011100000000000000101001000001000111011001101110100001000100000100110011111000001000011010011110101111111100010;
assign IM[16] = 1024'b1011000010100101110111110000111001110011010000011010101101111000011101111100010101110011101111010100111111000000101000101010001110000011011100100110001101111110111011010001111100111011000111110100011000011111111010001001001011010000011110100111100101101010100001100100101001001010000110001100110001010011010001010100000100001100010001001001000010011011111011010010111111101101000100000011001011111101010000111010001101001101111010001001111000011010110110011011100010100110000011011010000111101111001010001001001100011000111000101010111101100110110000010011100001100011010101110110011011011001001101011010000110000101111100111011010010101111110101110110100100111111010110110001001111011110101000011001001011100100011110111001101001011010100011101000010100101111110011001101110000000001101100100101000001100100100110010101010111001011101101101001000010001101110100011101010010110011011110001110000110001011100000100111110101100110001110111000101101111000100000111011010011101111100010001000010110001011000000011110010100100001;
assign IM[17] = 1024'b1101100001100000111111101011010000010111101011010011011010110010110111101001000000000100110100000011010101001111100001000001101111000011110111011001011111111001110010101001000011100100100010010110100101011000011100101001000010110100011100011000111010011110001000001010111111010111011010100100010010100010101100100011010011001000101110101111000000101101111011100101011100111101100100101101100110110111110101011011101000111011100010001011101000000001001111110011010010000100010110010101001001101100011001110010100110110100010111011110110000101100111111110001100000101100001010010001100101110111111110100000011110110011011110111001011010101000011001011010011000111000011101000010110010110001111011010111100100100010011001010001011001110111000010100000101001010111011111101100111100110111001001001010010001100101011101110110000011010111001100101000000100100010101111111100011100011110101000000001000010110001111101101101110001111011111000111001001111010011001010000100100110111100111110101000010110101101100100000010011000011100;
assign IM[18] = 1024'b1110110011111010011111001111010010000101101111100000101011110010101001101010000001111110101000110010011110001010000100001001100000000011011011011000111110001001110110001110001100001001111011110010110001011011010111001101101100100101011100000001001111011000110011101110100100101000010010101011101010101100011100010010011001101011011011000011111111010110011100110101011000101100011101100001011110010101010100000001000010100111111110111010110100001001000001110000110110101111011000100111101000100011110111101111010110111100000011011011111001111111001011001100110001000110110011010101010110110101100011001100100110011111101000000100001011100011010110000000111000111001000101101101000011000000000100100101001011111000000001010011010011000000111111010110100110100001111001010101011010101101001000000111111100110110101010010010000101011101001000000101110001010111111100000101110111110111111000101110100101111010111000101001110001001010010001111100101010111000000101111001110001001001010001001101011001010110110101100001011000111011;
assign IM[19] = 1024'b1011111101101010101010100110100001010110110000010110011100111000010000000011111000110010000111101100101101000010100001010111110000101110100100010011000110100000100011010000101101110111101000000101100011001110100001111110111111011110010001001111011101011111111111100001100001111111110101010001100000011100111100101101001001001111101010101111100100010011001000010100110111101001000011010010110001011100001101001111001111001110010011100011111000011011111010110001100101110110001011111100000100110001011011110111110011100001101001110010110010001100110010111111011000100101110010010000000001000010011001011000111010000101010011010101101001101000000100110010000000100110010010000001010011000101011101101100011000001001101110011000001101111100100110010010001111010101011010101010110110111110110110100111110101010101110010111000010000110100110010110100111011010101100001010101110001101011001100001001000010101010000101011100100011010111010001111111010100011100111010111000011101011001111110111111000100101110111101001001010100010000;
assign IM[20] = 1024'b0111111100110001101110101110000110110111011101111101010111111111000110101011101111010010111101000010111110100100110110101000011000101010011011100000100100010100001100011011000100101000100101110000010011101010011101110100110101111100110010010001101100010000110001111111100000011111010010011010011011000011010110111001101101010000111000001100111101000111010010100011000001000100110010100011111011110000000011011111110001000000010101001110011101111000110011010000101011010000101101111110100111110101110000001010011010011101100011100001111001011110010110011100100100111110111111011110000000110000101011100101111000100011110110001001011001100100110001101110100001110011110000011011111110100001011001000110011000011010000111100010001001101000110010101000110100001111000111111010101010001110100110010010011001110010111111111101110101110010010000001111000010101000000010011110000000100110110001101011011111000000110100100001010110000000111001111010100011111101100101010111000110010100101000000101011111110000010001100000101111010110;
assign IM[21] = 1024'b1110010111000101100000000111010011111110110110010001101100100011010110011100110011011100101101101110110110001110101110110111101110001101011011101110011110010100101010001001001100011010000101100000110010110110000000100110011101111110101000011100110000000010100101110001100011010011110001001110010100101111000001100001111010000010101101101111000001000100111100111100110111100110111110111111001011011111101100010101000000010101110010011011110010101101101101100000101011110011101000110101011011110001110010010001010000100001001001100011011001000000111100011110001101011000001000000101111010101011100011011001001000100011110001100011001001001001101110110101000100110011100110011111101100000000010000110001001101110100011111101000011001110001010010101001110110001101000001001111101001001100101001101110011110001111101111110101101101100110101011011101010111010001101010100010000010011110001010001110011011100000011010010111001100111000010001100010110001111110111000001111100001000110111000000110101000010101111100100101100111011001;
assign IM[22] = 1024'b0100101000110010111000111001010011010100011110001000111100110001000001100100110001000110000110101010010101101100101000101000011001001001011101011000110110011000000100100101001011110110000110110001110011100100001100010011110110001010000100011101010101110100000000000010100100010101000011010011001010100101100010001000101100000011101110101100001011110000101100011011101011010001010111111111000010110110110101000011010101101101111111010011010110011001110101010111110010101110100111100111111101111011011100001101001110010110000101010110111010011100001101100001101000010111101000000100101001010011011010110011000010110111011010010011111010110111110100101011001011111110101110111110110011110011101111100101000010010100000001100011100100001011111001011010111110011100001100011111100111010100001100010101000011101000110111010001111100111000101110011011001010111001000110100000001111001101111001101001110011100110001101001001101111001110101010101001001000001010101111100011010010111010001101111001001010000011101010101011001000111101;
assign IM[23] = 1024'b0010000101000111001000101101000011111001101011000010110100001101101111100111111100011011111101011000111001100010110010110010100010101111010011011110110011010011111110111101010001000101000100001110000010011111010000111011111110110000111100111101010110010001001010101111000101111010000000001101001011001101000001110110000100011100000101110111010011001010011011110010110001000001000110101000101010110110110000100001010011111000101101010011010110101010101011100000110000111111010110100101111100101100110111000101011001100110001011111100110101110111001101000011010000010001001000110000111100100110010110101011101110011111101011001110010100010010000000000111011000110111010111000101011110011010000100100101011000110111010111010110010111111001111101000100100101111010001010000100110111110110101100011010010001010011001010011110000101000100111011100000001010111101111010110100110110101111000011011111000011001000001110100111100000001010011100111010101011110101000000001011001001011000100110000100100111100011010110100111111110000000;
assign IM[24] = 1024'b0111100110100011101000001011111010100111111110110011010101101000011010000011011011101000000000000110000000011001011100101100100110001101001010100010010110101011111010111000100110100111111101101001110111110100000000001111001011101000010110010100111011001101111110101111100000101011001010101110011011010011000000111001011110010000101110111001000110110101110010010001101011110111101101100101110001100010101000111011100001110000111000000001101000000110100001010011101111010000010011100000011011110100111110110101000000100011100101001000101001100100100111111110111010111000001010111101000111111111001110110010110100001110001100101001001101011011110110000000101101011100110101000001100111101001111100110000010101111101001111101110111011010101000110100010010000100010001010001000101000101110100001100010001110011010100110101001110010011010100101010100000011001100011010001010001001011000101101001000011011111111101000011101111111100001101010010011110001000001011111110110011010010001011001011011111011010001111011001111110110100000;
assign IM[25] = 1024'b0010000001101000010100001110100100110000001011000110001001100001111001000100111011100000000110100111111001101110101011000111010010101001101100011100000111110110001100101000100110001000001101011101110010111000101000011011000001100101010010100001101010100000101110010100100111110110111101010110011101110111010001011100011100111010101011111001000101010010111001000000101100011011011000101011101100000111011000101111000011101000110111011100011010011011000001100001001101001010111110010011100010000111010000101000110011111000100001111001110110010010110010001011010010000111101000001011001011001111011110010101000010011111000010101010000100010010101011101111001100001001110011011111111011001101011110011000101000100100010010111101001110111111000100101011101010110011101111101010011000110001100000010100111100110110110001011111111100111110010101111101111001001000010101001110001010110101110001000011111100111100000111111110000011110000101110101101001111011101000111010100001010110101100011000100100001011010010110111101001111011110;
assign IM[26] = 1024'b0001101010010000000001011011101101011110011011000101110110101111111101011000100101011101101001011110011010110010111000101001000100101100000000101111110100101111100001011101011110101011000000010010100100011001000000000111011101000101100010010111011111111001001111100000001010100011011111011010111110001011001101101011101111010101110110010100100010001011111000111101100110000001101100111001000111100110001101000001011110011110000000100100010000011111010100111010110010011101000011110110010111010011101111110001010000000110011011001011100101101000000010100010011011001000010000111111010110100001100011110000110011110110010111000100101110111101101110001111000101000011100101010110110110111110101000010000100001011010000100111110001000101100001111011111000111110111101100100011111010000011001101010010010111111110111011100001100110100010000111110001011110000110110111100101001001101001000110100000111011110110101101000010011101011000010010001100010101110011001110011000000111110000101111001110000000011110100100011000110010000111;
assign IM[27] = 1024'b0001010010011001111110000110110100110000101011101110100110110010011000101001000110110101010001000110111001110010110001011001000001100101011100101100111110010001010011110101111100001111011110110111011010001111010101110011011010011011001111001000111001111111111011000001000101100111011000100011010001110110111011101111100100110001011000010011101001111010101001100110100001110011011100111001001110010111001011000001001101000011011110111110010010111011111010000110001000001110001100001100110011111000011101010011000001010111100001111110010101111011100100100101111011101111001011000000111010010000000011111111110111010100100111010101111100100100101011100001100100001010110001001001100101100010000011101101000000100010000011000100010101100100000111101000010010010100111111000011101001111110000100110010011000110001001001100101000010010110001000110001100110000101000110011100001011110101011011101011010001011000001001000000100111100111010111000110101010001110110101010100011111100100100000111110101001110001011010101111010011111011;
assign IM[28] = 1024'b0011000110101010010101000011000110000111110111000100101110110100010001011100110000000000101110001101110101001111010010111101010100000000111011111010111000111101111000001011101000101000101111010011111001110000011110100101101110111100000000001101100111001111110101111010000100100000110110100011010100110010000010011101011100100100001000000010000100111010001010101001011111101110010011001010010011101100111011111010000111001011101100110000111011000101101000001010001001111011100110101110001001011011011000101001010111100010010111110001100001000011100100001100011001010001111010101000010110111101010100011101001011000011011101011000101011110010010001010111110010011001011011011010101101001100010101001011001110101101110110000000010111101011001111100000011001101000011111010111100101111011011000111110111001010001000000100011101101110010100110110101001010110010000001011011001110001100011100100011000010010100011101001111101001111011011000101110101100111001000111111010100100001110110011011000010011111110100101111100001001011111;
assign IM[29] = 1024'b1011000001110010010010101000000010100011001101111111101001100110010110111010000010111010011100001101100001110110101000110001011111111100110010110110111011110000011010010001001100110100100000111111100000011111100111110011010010001011000111000110100011101000000001010111110101010001101010110000100110001011011101101110100101011100001101111101000111001001110011101100000001010010011111111001001101000010110100100101010100000111001110001110001101100000010011001110100100111110111101111010111100010101111110111000110100001011010111110011101000111011101011000010011101001011100011110110101001101111010011100000010011001011000100011100001000010010101000011000000000000001010011100100110111001101111100001110001010101011111100111011001011000101001101100101110100001001000010110110000101101001111111101111100110100011110000100101001000100000000001111001110110001110100001100100100011010101011111101101010111100010110010111110111101101110000100100110011110011101100001010001010000001010011010100001011111010110011101011111010001100001;
assign IM[30] = 1024'b0111111001111011000100011000010100011110000100001101011110011011011001010101000001111001001101001001111100110110000001110111010111100011010010001000110010011001110011101101010101010110010011110110011110000001010010110001011101000010111111010001011001111001001011001001101001111000100011011101100100100111111111011001101011011110100101011001101000000001010111011010111110010110001001000011111000111011100000100100011001010110111100111111100111101110101110000000110111000110100100010111110100000100010101110110110100000001100101111101110110110000010011011100000110001111010000110100100101011110000110101101101000011100111001011011110111010100001011001111101000010110110111010000000111110000100100111001101000111100111001111100010110010000101100100000011000001110000110101001111101001101111110010100100011111010001010110111110000110001100000100110000000101010000110101111001111101010111101101011100101100100010101001010001001000110010000111101111010011010010000100110001110101000001111111001110110001001001000110110001001100000;
assign IM[31] = 1024'b1011111001010111100111010100001101001110001110100001100101100001101001000100001001000000100100011001110001001100010110101111100101110000100011100001100111101101001110110010011010110011001111100110101111000010010110111000011100000011101110101110010111011111111111000001100000100110110100000000101000111011111011111100101110101111011010000100101111010110011011001001111111110011011100101000110111100011110011000001100011011011000101110001110000001110100011100001011110101110101010101101100101110100111101110000011101001000100110101110001000101010000011111101100011100000001100100000110111100111110110101101010111101101000100110000101000000000010001101010010000010101000111011101111000010111010101111101011100101110111010000111100000111111111010001101010101100001011101101010110110101101110100110010010111010110100101111100100111101011111010100000100010001100000100001100011111000100010001101110011110000010000101000100011010010000111101001000001011010101111010111101101110010000110100100100011000011010000111011000110010000100;
assign IM[32] = 1024'b0001101111100101000100001000001101110000010000110101000001110000000010000000101000101111011011011100011011110110110111111111011011100110001000001110111011101001001011010001011100010110101000111000010001101011101000100000001001011111110001001100110010100100110100100001010110000001110111010111100110001011111101001100100100001111101000011000111011011010100110100000110011111011101101100110100101110111001010001011100001000001001111001010101011001000111000101101100100000101001000110110111101011110011110101110000000010111111110010010111101101110001000101111010110000000010110000010011010011111010110111010000111101011001011011011101100111000111100011111011000010111011111010111110000000000000111110111000111100110110111100100100000110000001011010011101011100100110101000001011110011100010001011111011110100111101011111000100010000111101001001101001100011110110100100010000100001100011110000001000101110101011100010010100101000010010100101100011111101111111110100001111100110111011011011100001100000110000111001010110011110101;
assign IM[33] = 1024'b0111010001011001110110110011011011101011000010011001100111100010000011011000001010000001110000100010111000101100011010101011100111011010001011000110001111001001100011101001000010111000011011000000011110110101010010000011010111011111111101000110111010111110000111000010000010010111110101110001110001101010100010000111000011111010101101110100010000110101100101101100010111000001110110110000010001001010000001001100101101011010111001101101110111101100111111011011101100010101110001100010110010000010000100010111000001110100010011110011011100000110011101111010011001001110101001000000010110001000101000000000101010101111010010000101001110100010000000011110111010011110001111111111111010110000111110000100001010100110000101110010101110001111100011100111011011011010110100111000111101001111101110001100100100100011101101010111011110101111010111111001000101011011011011010010001011111110001111101000011010010010100101000001001101011001011011001001011110010101111000011110010100100010100111000011001111100100010111101111100111000000;
assign IM[34] = 1024'b1110001000000110000101001000010000100000011101101111111111001001001001110110011001010100111001110100101010111110111100110101110010110010001110001011100010101101101011100100011011000011011010001001110001110111010010011001110010000101001110101000110110001010011001001001011101100011110010111010111100101001000110111000100100111010100001001100010001101000111000110111111100110011010101000111111001011111111101010111000100011111010111100101010101101010100000111101000000111010011100100000001111110111111010101100100011010010011000001110011101011101111100110010011011010110100100000111010011101100100010100001010101011110101100100001011001011000110000111100001100101101001110000010001101010000011101001111001111011101111000101011001100100110001101001000000011010000011100010010010100110001101000101000111100011100100001100010001101110011001001101110000011101110110101010010011010010000101011000100101110001001111110100011110011001111001011100001110000101100100100001111000011000110010010101011111010111101111110100100111111101101;
assign IM[35] = 1024'b0111101000010100001000100101110000100110110000101010001100101000101001101010000101100000101110100100000110100010110110111110110111010110110011110100000111001100101000101011000011011101000111000011001010001111010111101010111000010000010010111110001101001101001011111100101101001100111001101100001001111010000000101001110101010111000101111000100011101001101101101011001110100001111001101100010001011001110010001111111011101000010100110110110101011110111011011101101111011110011110001110101011101111010011110011111011111010010001101101000011011000000001101111010111100011110011101101011001000011010111010111101100001111110011001000011001100011011001010011111100100000000000010101111010100001011101100111011001101101011010011000001001111001111000100110011011000011000001101001000011001001000000001100111001110101001100101111101001101011011101100001000101100111111010001011001000111001111101110100100010000010110011010000100011001111001001011000010101000101111000100110101010110000001010111101010001100000001010111010100001110101;
assign IM[36] = 1024'b1110011000111111001100011001001111111111010001110110010101111111101110010000001011011110001011111011111001101000011001111000010010011011100110111111110100101011100000110100001010100101010011101111001111000110100000110100011000011100010100110100000010111011100011011001000000110110010010000101000000011001101001011010011100101011111111000011010001110100011000010111101011101000110110011100110001111100011111000000110110010101001000100111001101100100110110001111001110001000000111101001101110100110011111111000010100001101001011100010111001111111000010111110110000010010011000011110100001111111000001111011011101010101001100001110001010011010010000101001000000100000111010010010001010000011000000110111111011001000001110111000011111100011001000101100011100010000101111000010001100010010010110100010110011000110111110101110011011100010010111111011100001010000110100110011101101100000011001111011001010100101111001110111001011001000001010111101111010001010100110010111001111100001000111110001011000110010001010101110100110101100;
assign IM[37] = 1024'b1010010101111101111001111010011111110001110001101011101101001011110000000101100000110101011100101001000100010101011110100001110011100001101110001001010011101001111010001101010010100111111110111110111000001100101011111000101010101000101011000000101110110101000110100010000100011000011010001111111101111000001000101001111111010111110111000011110001010101011010100011011100000110011010001011011110000101000100001010111010101101100010000101001110000010100100111010100001110011000101000101111110101100010110110010100011011010011001001111100011100101110110111110011100100000101000110100010110101000010111100101011010110100001101111101000110111111000001100000100101001100011000000101100001100000101101110010001011000100011100000101011001010010101001000010000110101001000110101111100111110010001101101011110011110111111011010111100101011010001101101100110010100010011100000100000111111100000000101100011101101011000101011101100101100011011000011010100110010110011111000101101011100111101000011111110110100100111000101101011001001001;
assign IM[38] = 1024'b0100000010101111001111011001011011011101110000010001110010010010000100001000100000111000111101111001111001110000000101110111111100101110111111001010011001001111011110101110011011111000001011001000101100010111000110010000110011111011000001100000100001011111110001000110001001011011110110001010100110111011111100111110100000100001111100010011010011001100011011000111100011010111001100101101001011101110101000010011001111010100011101011111111000110011011011111110100010110111010011000010010110011100011001000111110111010001011000111110101001111110100001001001100011100010000001000010111001000101101110010100000010010111101111101001111110010000111010010111011100110110001100001000000011101001000110011000101011000101011000001011010000100101001011000101010110001010001100101110111001000000000000111101000010110010111101100001000000011010001011011100101101001110000110010000110000011111110111101101111111010000011110110110010011111010110110110010100000000000001111010010001000101010110100000110011100101110111001101111110111011111;
assign IM[39] = 1024'b0000101001101111011001101101001100010110110100101000101100010101000111111011110111001001101110111101101101000001110101001110101110001011111110001000110100110010101010001110000101110000011010000001001111011110010010111110010001110101010100001000100010001110010011100001110110100101011011011101001110011010011110111101010001101100001100100010110100001001101100001111111100001101111011111010110011010100101110001000101000000011100110010011110101010110010101111100110101001000101000000101110100111011010110000101111011110001010110101001011001111011100111011100000101100100100000101001011111110110011110001000011100000111100111000100101000000000011011000101111110100011111011011111101100000101011100011100001000100101000011100101010010010100010011000010011101111101001110011100000010101001100010110100001111001110001010011100110000111001010010000001010100110101001101010111110010111000000011111110001101101111010001101100011000000110101001111000110100001100100010101111001101111101110000010010011110010101111100010000110001110111;
assign IM[40] = 1024'b0000011000101000110000010000010110110011100010101110001010110001000100011100011100100010010111011111011100101111111010011001010001111101011000010110101010111101001010001011001110001000001111111111110111110100100100101100001110101111001000101001110001010100101100010000010111101101000001111000111101001011011010110111010000111101111011101001111100011110010010110010000110001010110100110101010101110001111101010011111001101011010110011100001001000001001110000000111011000011111000000100011111001110010110011001001101011111111010010100011001001101110111001110101101010010000001010101100111011110100100011000101100111100101011100111110101011111100001011110010011001100010000001000001111101000100110011000100001011100101110101001110111100001101110000111110010110100100001001000110001000001000100011100011101101000001010001101110101011011011010110011110000111111000001110011000111110111000000011000000101000001001011010000111110111111010010000011101100000110011101110110101010101111111001010011101100101100110000010000101110111000;
assign IM[41] = 1024'b1000110100010101111100010101110100010101000011000010110001001011101001100111011001101110000101101011011101011110000000100010110011001110111001111010110011100100111011001011011000001100101111000011111001111011011010000001100001111100100111110001111111011001111000010011001100101000111100000000010111011111011110011101011001111111111011001110001110111000100111000000011010010011110111001010110110011100111010010100111110000100010111110010111001011100010110010001100001011001010011100010001100010110111000010101110000101111000000110011010011101010011111100100010001011010110001010100010111001111101011001001011011100000001011010101110110001000110110110010011000011011110001110000100110100010011110110000111000001010000100001101100111101000100111010001011110010001111111110100101001000110010101010000011001111001110100000010100011010000010010100010100011110110011001010001101100010111000000010110101111111011001000000001001100010100000110000110111100101001011111101111001111001100110011111110000000101101111100000101101111000101;
assign IM[42] = 1024'b1011000000110110101111100011001110000011001011001010001011000001101001001010110010110111000110100000001010010001011000111000100011011110101100010011101101110111010010111111001111110001011111000100010110111011000011111010110011110011101010001000000010101001000010001110001011010110011110111111101100101100010110001011101010001110101011000000110001100111101010001110101001000001110111100011100110000100111000000101101110110110100111001110100100101010011000000000001111010100000111111100001101010001011111001001010010111110110101001011001111111011010110001011100111001101111010001100001111111101000110101100111010010000110101001011111111111011011100001100010111100101011100110000010000100010101010000010101111110000100110010101010101001110100100101101000000100000101100001010110100110010010100000101100110101011100100100011111011111000100110110001111110111100101111111100100001111000101000001111111000000101000010110000101010101000001000011100100011000110111101101000001100111011100101100100001001110001111110001100111010111111;
assign IM[43] = 1024'b0101100110111000011100011110001101011100001010110111010011100000010101010001111111010111000100101111110011110010100101001101010100101011111011011101001000001011111000001100101001111001001101100010110101110110010111111011110001000000111100001010000000110011001001010110011110101101011111001000100101110111000111000100100010010011000011111011011111001101101100101101001111001011011100111010100011010001111001101111001110100100111100001001011101000011000100011010011111100011010011001011011000000000010110010110110101000111011100100101010100011000011011110101100001000001101110001111101010000011010010011110011001011010101000000110010110110010011111111010100010101111101111000110000011000011001001010010000001010010000000110101001010000010111110000111111100101101011110011010010101011100010110001100110100110011011110001010110011010100111101101110011001001101010001001000101100100001001100101110010001001111010111110110101010000000101010000010001011000011100011001101111001000111111010011110011011011111110000000110010001000111;
assign IM[44] = 1024'b1001001000011101000000010100000011111010110011001000111100000000000011010110111010010111111101011101010111111001110001111110001111011000000000100111011010011101100000010110011111000101000001000010110000111110001100010011100011111100101111001100010101001001011110011000100111111000000001001100001001000100010100011011111101001101110000111010101100000011000010101110011011101000010110000011000111011010011011001101111111101100111001111010000100110001101000110101010111011011000011101010111110011010001001001001111000011010011100111101110011100011000010000110101100010110100111011010000011010110000110101100000010001110010001100101111111001100000110000010000000110101111101011011010110101110110011000100000101001110011000111010000011000001000101010111110010011111110001000111011101000101100100010101000111101000100101111100101010011111010101110001111010100110110011110110110011110111110011111001100000100011110100010101110100011000111101010011000011000111111011111011001011101011011000100001101000001111011100101101101111101000;
assign IM[45] = 1024'b0101001101001001011101101111100110010011010111100111011101101010010010110101100101000001110111110110011011001110101010101010101111011111000110011000101100100100001111111010011011000000000100111011100111110100011011110001101011101111000101111011100011000001010101011000010101100101001011110111000010111110000101001111101010000111011010101010000111001010011101000100110011011010110101110000011101001100011100010001010000010101110100101000100011000000111100010011101100111000101011010010011100010111110111100010101000011100100000000110010110111101010100011000000010010001111011000100011010101011110111000010011100010001101001110000110001010011100100101001011010000010100101110000010100110111010001010101110101111111000100110111011010101110110101001101110100000001000111111011111001110100111110001110011100000000100111110010010000100011000000111011110111001000101100101001110001100001111111110111111110110101101011001101011000011110111010000011010100000001001110100011001111111010000000000101000111100010001010001111100000011100;
assign IM[46] = 1024'b1010101000011101100010111001010101010011110101110001101001100001100000010101011000011100000110001000001111011010011110001101001101100011001101001010110000000110010000110101111111111011011101100111000110100111011000111010110000011011000100011010100100101110001001011010111011100000001111000111100010001101111100100110001000001110000101101010000011101100001111011000011011111110101110110101011101111000010100011001000001111010000110010100100010001011100011100111101110101111011010110100001110000101101111000011000001111011000100110000100110001010101001011100101110101000110000100011110010111010000011110000111001001110001010010111101100111011011101110001011101111000011000001010101000100101001110110001110111100000010000001111101110011001110100100001111001110110011001010110101110111111010011101010000110010000110001100110001010000111011001101101110110101011000101000011110101100110001100111111100111100000001000101011010001111110011001011000010100110011111010000111111111111001100010110100101000100111000111000100111010101010;
assign IM[47] = 1024'b1001001011000110111001100111100010000010000101100101010001011101111001000110010001010110000100101110010001000101101110111011110000111010001101100000110001010010000001111001001100101101111111111101000011100011010000111000001110001011000011011000100001011101011000101001000000100011110110000001000000100011101001101100110010001010101010011000011100011111111011010101101111110000011010001000010000111001000001110101011101011110010000000100010100010001011010110101111110111000100100001000010011001011011101101001011100001100101110000101011000001011000100010100011110101000011101100111101001011110001111111000111101010000101111101101011000110111110011111011101001000111110011111100100100111000111001001110110011101101001111100110110000110100101011100000100000010110010101101001110011111100011011000011011110111011011111111110110011010111001111010101101001100110110101101100111000001110001110011110100101100000001010011001011101000110110101001101111111101010000011001111110110010101110001011010001011011110000001010101000000011110;
assign IM[48] = 1024'b0110011111010101101111111100110101010011011010110101100000111100010011110111100011011101010000000000111111000101000111100000111111010100011111111011101010001100011011010111111111110011101101100001010001101110010010101110011010111111101000011100011100000010011000011010110101011101010011111110010100100110000110000111001001100010110001011001000110011000010001010011000010001000001010001001110101100010001001010010101110100110011010010010110111111111101100111110010110101101111000010100010111010000011001101000010101101001011001101010101001101001000010100101011001111001100110100101100010100001110100011111111011000000110110010100010000111111000110001000000011100101011010101111110011010110100000010001011101110000111111011110000110001001010011110010011110011110001110110011010000100111001001000000111101110110111101101111011001000111001000000100001100100011010111100001111010110001100111000100011011000010100110111100011100111101100101001000100101101100110000111111111101000100011010010001100001110000001001010000110000100011;
assign IM[49] = 1024'b1011011111101010001010100011100100111110100000010011100110011011011001101110110000010101001111000111100011101001011100011100000111100101110011001000011010001011110000100001010100110010110111010011110101100100001100110101100110000001001101000000110100011110110011011000101011000010011111100000111111000110111110100110100001100010101110101000101001101110111111101001010100001010100111000110000010100011011001111101000001110111100010101001110100001110110100111000011001111101000100010101110111100110011111001111111001011110100101111001111000111101111111100011010101001000000110010010000110101011011010000100000110001101010001111010000011100010010111010101101100001000110011011000100110111001011010000001100100100100100010110101010010111100001001001110101011101000100110111110101000101000111000110100111100011101010101111011001000010001100001000111101101111011100110101100001001000101000011000100110011111001100110011010111101101000100010101001001010011110111101101110000011100101100101110011000100010101001111101110011000011100;
assign IM[50] = 1024'b1010100010101011100101010000000111011001101101001010010001001111111001100000001010001010010001110000000001101001001011001110111111010111011000111101001110010010010101010010111100010111001101001000001111011010010110110000010111011000111101111100101101001100001011001000101111111000100100101101101111100010011110001001000010010100111100101001100110010110000111111110001101100101110010000110000010101000110010010010000011111001011011010010111111110111000011001111110100011111010001111100101011011111011100000110111001110000011111000010010111111010001100110101000011011011001101011100100110110011110000010001001101110111101011100111000001110101000100011110001100010101110001110100100111011001001001111010101001101110000100011000101101010101001010100011110111101010000010011000111001111000101001110000100101110011110001111111100101101010100000001100110000111110000110011001111000101001010100101001110010110011001001111101000011111000011000000010000101000111100111010101100011001101110110110010011011011100010001100000111010001011;
assign IM[51] = 1024'b0000111101110010110011000110110000101111000110100100010111011011010111011101101010011001011011001101011011101100011010001011011000010001100101000001011110001011100101010011111111011111111001001011101110101010000000001010110000110100100010100111010001001000111001011001000111010000111000101110000001001100100101100111010110110100100110100100001110001000001100001111111100001001010000100100101110011111011001010000101011010010100011110011000101101011111010100101101110011011101001110100111001101100011010000010110101111001000110011101100011011110100110011110011010111111110111111001010010001010011000011000101011011010010100001100100110010101011011010101000011000100110100011011111001010101101100100010110011011111001001011110111111101010111001110011011111001000100011111110001110110011010100000001001100001010111010100011101000111010100011000110010011000011000100111000101101100011111101000011000001000011101111100000000100011011101010101000110100100010010011110001001110000111100111100010100010101001111111001100110100001001;
assign IM[52] = 1024'b0111001101001000010001111111111110101111001101101111100100011101011110001011110110100010001010000100111010001110111111100001001011001101100101100001001011111001011010100010011100011010011100010101110111000110010011011111000100111111000011111111001100011111110110000000000010111100101111101101001011001110111101111000000101100011000101101100001101011111010101010101011110100111100010000001000100000001001100100010001101000100000010001011011111111000010101111111101000001111101100111101011101111001101111011011011010011010110001111111100011000110100001011010001100000000101100110001011001110001010001001110000011000001011000011101001110111111011001010010100110110110010100110000011010001100011101000100001100101100011101101010110000101001101000111000000101110000111110101110010101101000111101110100000010110000000001101110100000000001001010011000001101011100010001101101001111111011001100111001010001100101100100000100000001100110111001100011010111011111111101000011011101010000100110000010010000101111011001001100110101011111;
assign IM[53] = 1024'b0001111111010001001011000000111000100010100111101001110100101110010000011101000111111011101000110000010010101110111101100101111011111000001000000000010101001101000110011110100001101001001100011110000011111111010111010000001011011011011111001011110011100001100100001011111101011000110111001111011010111011000001010100100100111000010100010010111101111011110010010101100111010111010001101000001111001010011000001111101000000110101000001010100100110110001010100111011011011101111100111110000011000001111110000001101011000101001110101010101000111110100101100100110100110000001011100100111000001111101010010011111001000101010010100100011111111110000010010000110110011101000011100011000010110001110001100010000001001011100001010001110110001101011100111101100110001101110100000001110010001101011101110111000011000110111111011001100100111000010101010010110101110101100101111011010011110100101011111101010100111101000111011101100010001000100100001010000000001111101101100000110101000100011111101100001100111100000011111011100111111001;
assign IM[54] = 1024'b1010000111001110111100001011000111010100011011111010111110000011010000010011000101001001010100001001111100001100100010100100000111111100011001001100001010110001011111011110111000110101111110100011110111100100010010011001010010100100111011111010000010000010010010100100001000100001101111011100001000011001101101111001101001000011000011101100100010110111011101111101011001100001101011100001101100110010110010001111110100010101001101001000011010000100111011010000111100110010011111000011100010000101100111111110111111001100111011100001111000011101000000010011011001100100010000110001011110001111111110010001110111001001000010010101001101101001010110010000001101111101011010101000000000011010100101111010001001101100011101010011000001000001010110111100111111111010001011111111111111111100111100010110111010010000010100100110110111101000101111101001010011111101100111100001010000000110010100110101010000100001001010110010101100101101110100000110111011001010110111001100010100000100101100001111100001111011111110001010011011100101;
assign IM[55] = 1024'b0101011010011100001100001110000101100010110001011011110111001010111010110011111010001011110000111100110001101111000111000110000111101110011010100100101010011011100011010011011110010011101011100111010011000100011100010101110100110011000110110111111011101001110010001101110010111011110000001011011011100000110010110101111100100010100001101010110100010011001010110110010010111101100001001010110110110111011110010011111001000100000011000110011101101111101010001001000010110001110100011110101000001100110001101110000011000111111011111011010101101010010011101100110010000111100001001000001000101100001010010101000000110110111000100111010110000101101101001001101111010110100010000100110010010000000101010010010001101110111011110010110010011001111001101101001000110001111110100010011111110101100000001001111100011110000010110011010010000010110100110111000010100110111000111011111101000001100110111101100010110110110100010110010000001111010001010111101010111101101001110000101000100100111011111101000001100000001001011010001000010111;
assign IM[56] = 1024'b0110000100110101010101011001111110011111011011010100101001101110110100111110101101111010000001100000101010101101111101001111110001001001100111000100001001100101111001111101110000100001101111100101111101101100010000000101000011101101110001010110001001001001101001111000111001111001000101110111100011010010010110001011101000101000000100101011011011101111000010000010010000110110101110100111010101010010011000101110100011001011101110010101100000010110010011100110110110100011000101110111100011100100110100101101011011101101001011000000011001110001110101001100111000011111011100011100100101100101001100001010010100000100001111101010100010110101111010100101000111011011011101100011100100100000101111001100010000010110110010010011100110111100011010000010111010001110001010100101110110100001111010000011111101110101011100100001011010010110010100000110011100111000000100101110100001101010110011101001011101111111110010101100000100000110110001011101111100011010110001110010001100000100111110000001110101100001011111101101101100100010;
assign IM[57] = 1024'b0111011110001100111101111111001100011111001001010010110001001100011110100000110111111000011110110101111101100111010111010111101101111000011011100111011100000100111001000101001110011000101010011000110000101100100110111011101110001010011100010010110001011010001000100111100011100011001111010110001001110110110101000010010010001111110101111110000000101101111000000011111101000110100001011111111010001010111101000001101110110100111010011101101010011000110001100101111001100011000111010010000111101110100001011001011100001000101000100101101000111011010100010010011101001101100111110101010010011010010100010001011110110101010110011001001110011010000111001011010000011100011100000000110100001110010000010010101101111100100011011110110101111011100100101101011001000101110111000100001000000110000010110100010010100100000100000010011110100001000100111100100000001000001001101000010111000111111000101000100010101100110111010100110000011001101100110111111101111011001111001010001100110001001111001100111011101110010100111010110101110101;
assign IM[58] = 1024'b1011110100101110001100010101001110000101111100100110100001011110010010101001010001011100111111100111100110100101110011001110100100101000011111001101000110001101111000001110100010001101100110000111001011111001001011100110010111000111101010101110010100000101101001011011101011111011101000000100001110011000100001000000101100000010001010011111011011011100010101100010101001110100001011100111000011011101000000000000111010011010001101101001011011100011011101011010001010110011110001000010001001000111110011101100001101011101000111101010001100100101110111110000111001110101001111111111111000011110111001001111000110111111101100011100010011110110000011111110000001010011101010100110010100100011111000000010110010110010111111001111101010100100111111011111001110010000110001000110011110001010000111110000000000110100000000111001100011101111011000001011111101100011011110101010000001000001010101101010011001111010000101101000011101110010010010001110101110010111011010101000101000110110001111111101010101100101010000001101000000100011;
assign IM[59] = 1024'b0010010010011010100001101111111101001101101000010110011010010010001011100011010001010100011110011111000011111111011111011110100010100000001010110110011011101011110001010111010100001101011101100000010111100101011001000100000000010000100011101000111111010001101000101011010010100101011010101110110000001011110101011110100000001011110000110100110100010010101111000001000000111111100010111100101101010111101011101001000000111111110100101001111010011000101010101010011010000011000011110110000110111111101000111010111010011101100111010101100001100100111100100000010000110101000100010100110000101111000010011100100101001010101111100000101000010101000010010100100011110010100011010100011101011101100110011111000110001111010111100011100010010000101110110001001100010101101000010001011010010001010100011010001111011000111100111111111001111000000111010010010110111000010110111011110101110101110100000110101000100000101011010110011000001011011000100111110100011001101100011110110110111101010001100101110011000110110110111111101111111001;
assign IM[60] = 1024'b1110111100101001100000110101110101110011000111100111101110000011111001101100100011001011010101011101000110010100111100000001101101100101001111111011110101001110101001111001000111101101110101010010011100101101010000001011100001000010101100100000000000111011010111000100010000011000110001011000010010100110011000100001111010110010010111100100000101000001110111000100000101001110101101111111010100111001001101110001010010100111101100110000101010011010100000111010000010101110001010011110001011100001101110100001000011001101010001011000111111001001011111001101110000111001000010010000110111111101110110110101010110000000110110111100010100100110101001010100100101011100111010101010011101001101000000011000101110101000110011111011101011111001110100000100010110100111111110001100001011000101000000010010111000110000111110001101100011110011111110010110001010000111101111110001001000101011111011101111110111101111110110111010011110011110110110110001000101110101000001000000011101001000001010011000011011100100000101111101110101110000;
assign IM[61] = 1024'b1111001100110111010110000010110000000101001000011011101001011110100110011000110001101001011101011100110101111111000101010010111101110010000010100010011000101100110011100010011001101101011001101110011000000000110011011011011011000100101111110000110110001001000001000111010111010100100110100100000001110000101001010100001011101001111101101001010101010011101000001101000111100000001100010011000011101101011100100110001110001011111110010110000110100110100010100010011111000100000000010001100001111010011000110110101100110000000100111001010010101110000010111101110010010110001110010011110001010011011111000000000001010001001110001011111111011010101101111110010010011001100010011000100110100111100001011100110111011101101001011000110111110100001100100111011111111100101010011001110101111111111010101000110101110100100111111110001000101001110100100110010011010000100110000111010000100001110010110110001100000011110111111111000011110110100111010111111111011111101111111001011011100110001001001001100010011010011110010000101100010100;
assign IM[62] = 1024'b1111110010111101001001010010101000100111000111100111000010010101001001111110010101001111010010011100000100100011010111011101001001010111010001000000000000100111100000000011011100011110000101000010111100110100111101001001010001000101010111000011110101010110010000101011110000011101001100111011111110110101000001111100000110111000010110100101011110100011100100010011001110100011111101000011000010001110110010010101100000101011001110011100000101001011110100110110000101010010111010101101101001001001111110010111001101110011001000001010111111101100100111110010000101000010111011010110010110111011011101111110001001001001100010110101101000101011111000011110011100111001110001101000111100011010110100110101100011100101110000001011010111101111110100110000011101111000001110100001001001111111110110000100011000000011101101101110111100111110010011011101001000110010010111110011101010111101011101011000100100010000101100110100001010101000110011010100010100001010110101000110011101000110000001111010100000110001001100011011100110101111;
assign IM[63] = 1024'b1001010011110110111011101100111110001100010011111001011011000101111001101101110000111011001101010110010011011001101010011010000010000011001101100000110101101011100001100001001001100001100001101010000010100110001001100110111100001000011000110000011110001101100010001010110001011110101011101001011111010100100000001101010100101110000111011011001111111110110001011011011110100100111011010001010011000010001100101001100000011001011101011010110100000110101100111011100101101001000001010010110001110010100100110101001100000111110100000111101011110001101110011000110001111110110100010010011000011101000100111001011101101100101010100111111001101110101011000111011101010101000010000101000010010111111001101101111010000101000111011001100000100110011101001100011001000111110100010010011010110001001101101110110110101011000001001101100101010110001111010101110111001100010010111011100010111111000011001000100101010101101011011000110101101000000100101101001101001001111000111100110101000010000010101110111111001100001111111110011001000111;


//LUT
integer i,i_cf,j;
always_comb begin
for (i=0;i<E;i=i+1) begin
    case(LBP_codes[i])
        'd0 : LBP_hvs[i] = IM[0];
	'd1 : LBP_hvs[i] = IM[1];
	'd2 : LBP_hvs[i] = IM[2];
	'd3 : LBP_hvs[i] = IM[3];
	'd4 : LBP_hvs[i] = IM[4];
	'd5 : LBP_hvs[i] = IM[5];
	'd6 : LBP_hvs[i] = IM[6];
	'd7 : LBP_hvs[i] = IM[7];
	'd8 : LBP_hvs[i] = IM[8];
	'd9 : LBP_hvs[i] = IM[9];
	'd10: LBP_hvs[i] = IM[10];
	'd11: LBP_hvs[i] = IM[11];
	'd12: LBP_hvs[i] = IM[12];
	'd13: LBP_hvs[i] = IM[13];
	'd14: LBP_hvs[i] = IM[14];
	'd15: LBP_hvs[i] = IM[15];
	'd16: LBP_hvs[i] = IM[16];
	'd17: LBP_hvs[i] = IM[17];
	'd18: LBP_hvs[i] = IM[18];
	'd19: LBP_hvs[i] = IM[19];
	'd20: LBP_hvs[i] = IM[20];
	'd21: LBP_hvs[i] = IM[21];
	'd22: LBP_hvs[i] = IM[22];
	'd23: LBP_hvs[i] = IM[23];
	'd24: LBP_hvs[i] = IM[24];
	'd25: LBP_hvs[i] = IM[25];
	'd26: LBP_hvs[i] = IM[26];
	'd27: LBP_hvs[i] = IM[27];
	'd28: LBP_hvs[i] = IM[28];
	'd29: LBP_hvs[i] = IM[29];
	'd30: LBP_hvs[i] = IM[30];
	'd31: LBP_hvs[i] = IM[31];
	'd32: LBP_hvs[i] = IM[32];
	'd33: LBP_hvs[i] = IM[33];
	'd34: LBP_hvs[i] = IM[34];
	'd35: LBP_hvs[i] = IM[35];
	'd36: LBP_hvs[i] = IM[36];
	'd37: LBP_hvs[i] = IM[37];
	'd38: LBP_hvs[i] = IM[38];
	'd39: LBP_hvs[i] = IM[39];
	'd40: LBP_hvs[i] = IM[40];
	'd41: LBP_hvs[i] = IM[41];
	'd42: LBP_hvs[i] = IM[42];
	'd43: LBP_hvs[i] = IM[43];
	'd44: LBP_hvs[i] = IM[44];
	'd45: LBP_hvs[i] = IM[45];
	'd46: LBP_hvs[i] = IM[46];
	'd47: LBP_hvs[i] = IM[47];
	'd48: LBP_hvs[i] = IM[48];
	'd49: LBP_hvs[i] = IM[49];
	'd50: LBP_hvs[i] = IM[50];
	'd51: LBP_hvs[i] = IM[51];
	'd52: LBP_hvs[i] = IM[52];
	'd53: LBP_hvs[i] = IM[53];
	'd54: LBP_hvs[i] = IM[54];
	'd55: LBP_hvs[i] = IM[55];
	'd56: LBP_hvs[i] = IM[56];
	'd57: LBP_hvs[i] = IM[57];
	'd58: LBP_hvs[i] = IM[58];
	'd59: LBP_hvs[i] = IM[59];
	'd60: LBP_hvs[i] = IM[60];
	'd61: LBP_hvs[i] = IM[61];
	'd62: LBP_hvs[i] = IM[62];
	'd63: LBP_hvs[i] = IM[63];
    endcase
  end
end


endmodule

module BINDING # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  [E-1:0][D-1:0] LBP_hvs,
    output [E-1:0][0:D-1] bind_outputs

);


logic [E-1:0][0:D-1] EM;

assign EM[0] = 1024'b1011110011000000010100011001100110001100000111011100001110101001001111000101101110001000110110111100100110000001101101110100010111110111100100010001001100000101101001101000000001101001000100010011011010010011000110110110011010110000101000011100111001011010100010000110100001011110000011111001000000001010100010001011001010001100110111011100010001100010101001111011011100000011110101110000101010101001001000010111111010111100100110101110111011011000001010000101101001100100010011000010101101010100011010001110101100101011011000101011100000111111110010100111000000111101010000110101110000010011010110111000111110111011011011111100011100000100100110010100101000100101000101001011101101011011111000101110111110111110011001110111001101111001000110011111000100010001000001110101000010110111101101110011000000001110111000000111110001111010100110110001101101101000100111001010001011101011110101011011001001100010100001111111101001101000001100101010001111011010001001111101110110110011101110011111111111110000101110010011100111001101;
assign EM[1] = 1024'b0011010110110111010101001111010001001000110111001000110100101110100100011011100001011010011111111100101011110010001011000010101111110111000101100000100000100010000010101001100011000111110110011001011010010100010111101101001101110110110111010010101001111011111110110111100101101101100110110111111111010100100101111100110100011101011011010111010001000111100011110011100110100101100010100101101100011011111100101010000001100010011010000001101111010001110001100011011101111100011001111101101000110000011111010100100110010100010001001000110111010010100110010010011110010010001101001100100010000010010101000011100001010101011010001001010010010100000100100000100101000000110001001011011101011110011110010100111011001010010111010011010000111111010111010101111011010111000010111100101111011000001000110001110011000110100111100101100101111110011010001000011110100000001001011000111010011110011111100000011101100000010100110100110010011010001010011100100111010101010110111100000100110111101111001000110100000010000000001101111001001111;
assign EM[2] = 1024'b1100110101001100000000101110101110110110000011100110000100101001111001000100101110001110001000011001001000011101001100100011011100100111011001101111000111010100101100100001111100100100101111101011000110110110101000100100101011101110110010011110110010100111111011100001000010110010010001100001101111110110111111010100101101010111110110011000100001001100100101000001001110111010000001010111100111100111101100010000110000001110001001011101111110100110101000001111001011011010000010001110111010110100011011110000110011110010011010001010101111011100111111001100001111111001100000011111111001110000100101110001000101001101101000110001111111001110011000101100001001110110000001001000111100001000101011000010011000010110110100100111000110001011101000111010001110001011011100001110001010101000111001001011110011110100110110100011101001101001100111001011101111000101011101101111010010000101111101100111110010101100000110001110100001100011110101111001111000100000001100100011000001011001010111100110110001100010100001101100111011100001;
assign EM[3] = 1024'b1100000100110101010110110110011000111011000101011000111011111000000010001010010100110100100111110001111010100010000011110010010110110010001011001100011110011010101100101000000011001101000101001100010011011111010111010111000000110001000111110110010000000110100111111101000001000001001111101000101010101011011110100010000010110010001100011001111110010011110101110010011111001101100111001101000000011011100011010011101100111001011110000110101101000011011010000110111110101100100001011010100001100101101100001011000100111110100000111111100011110111011111110010111111001100011111100010011100000111111111110010010001111000010100110010111000010100100001100011111001110100110101111000111000110011111100111000100011011000010111010101000001011001000010011111100011100001100000101100100000001100010111010111100000001010101000011011111101001101011001111001110011111100010001001100001111011110100111110110101100001101000101001010101010110000011001111100000001000101110001111001111011101000101011001010110010111110010110110000101010111000;
assign EM[4] = 1024'b0011100010010001001011111111110001100101010011100011110011001001010000101010110001111001011101100001101001101101101110010001111100011010011011111011010010110001000011111000011001010111010011110000001000011111100110111101000101100000111010011111101110110100001001100000001000010001011101110111101111010100000100110101100111010101100000000001101000110011101011011010010001100100011110111100111011110101110000101000000101110011111001110001100100101001000111001011111100111100100110000110000010000001110001100001000001000111110111011111001111110100101010000010000110100000101010010001010100101010101000100010001010111000101100101011110101000011000101011001110101001001010100100101010000100011101011011011010011101001100100101111001011000110000111111001100011000001001000111010010100110100110011100110010001111011111101001101001111111000010110000111100100001011010011110001010011011010111111011111110010101111011111011010001001110000101100000011100001111101111111101001111100001101010010011101010100100001001001001011011000111110;
assign EM[5] = 1024'b0101001000010110111000100110011101001111100101000011011111001100000000010011101011000001101111110100111010011101001001000000000111001011101100100100110101011010110010110101000100011011111100001101011010010001001011111111110110101110110000111000010001001000001100000001101011111000110010101101101011011110111010000001110101111110100100011001101101010101011000000110010101001010011011010000111110101011010011101011101101100111100001111111100100001011001101100011111100111000001000111011001111100011110100010101011100000110110001111011110111011011000010001110101010100101001001001011000100011101100101001111101011010000001101010010100000111011001010101000100111101010011101000100010111100111101010100111111100000010111000100011001001011000111001000010001010110100100001110001111101100100110110000000010100111111000000000100010111001111100110001111011010111010011110111100110011110011100000101101100110101001011011000000011111010101001101000101011111011000101010010010111100111111010000101100100000110001111111001101001001000000;
assign EM[6] = 1024'b1001010111010100000000111001100000100111101100111101000010101110110010100110011101011010000110011101111011100101111001000010011010111101000100001010111011010100100001111111101011111101110011011001101001001001001111001000001010010001100110001100111100011111010000001001100100100010001110000011101000010101110011110111111100010001000110111001101100010100111111100010111010001111011110011001101110111101000110010000110110101000111000000101001010010110001111010111101001000011101111110010110111011101110001011011110111001110000011100110000000011111111110111001001011110101011011010010111010101011110000001101001110010111010101011001001101101010101000000101011101110011001101101010001010111011011011111010011101101001101000111110010101111110111010010001010001100000001100101100100000111111000111010101001110001101101000000001100101000100000011001101100100001010000001100001011110010111100000001111100110001100100001110101001110001101001000000101111000000111010110010001001000110110001000100110011111100000110100000000011111101100;
assign EM[7] = 1024'b1111010010011001000010001101011100101111100110010000101100001010011011000110110001010000110011111011101100100111101110010010001011100000110000101100111001111010111101101001101001110011101011010010011001001110011001001001100010110000100011100101010100110110001101010001100110001000010110100100100000001101010101001001001100001100001100101001100001111111100110010100100111011111011101100110111011111100000110101001001110100101001101001001000110010100010010100111011101110001100010011010110111110110110011000011100001000101100110000010110101011111011011110100010010100000100000101010011010111011101000110001100110000010101101010111100100101111010110000100110000101101010110100001101101111000110110010011011101110011001010111011111011101110011010000011000010110001010010010111000110000000110000110001001011001101001011100000110011101000111000001011110011011000010001111110101111110101100110100101011010011111001101101100100001001011111111010110111100100000001011111011110001010010100010111001101110010101011101111001101100011011;
assign EM[8] = 1024'b0111110001111100001101100110000001111101001011110000011100100101011001110000011100100001010001001111100000010000110111110111001010000100111110111111001110111110010100010110001000011111101010001010101100010100111010110111100111100111100010011111100010111101111111110000011100011000111111011111100001001100111001000001110101011100111110011101110110010101011010110001101100100111111000011001000100101001101100101110100001110011011101001011000100001011110000100001100101001010010001110011010111101001000010101011001011111001100010000101010000101010110010110101100100010010101010001010100101000101001001100101001111100011011011111010000101001001111000000011100001111011011101000100101100000100000111111010110110111001111110100010010001010011001011000101010110000111000010101010110111000001100110010010010011011110111010000100101111010001100010000011000100011110010101110000100100001011010010011000010010111010001010001101010111001111111011101000010110101110011111010011001010010001100111001110011000111111101010000001100100111110;
assign EM[9] = 1024'b0100001110101010001100011001011100110100110110010100111000010100110001001001111001100001011111101000010001010111001010011011110110001001011011010101011010011110101011101000111100101001111100010000010111111001101001011001101011010111100111011010110000011001100101101001000111001001000110010010000010100010101011010000011001011011000111010010010000000001100110000111011000110111101000001011001010000000100010101100101101110010111000000011101110010011101011101001111100011110101100101011111110001001111101001000011001010001100001101100000101100110001100000101111101001111100001101010001101000101110001000100011110100000110011001011011111101100111111000110010001111011100100000110010000100011010111010000101111110001011000100100011101101010000110100011010010110011011110011011010100001001010100101111011100110000011010110111111101011000111010111011100010010101111100100100000101010011011100110110111011111101111111100001110010101110111111100010010001101101110001101010100111110010001101010110110000111101011010110000010000001011;
assign EM[10] = 1024'b0111001100111110011101001101110111001010101000000111111010111001001001111100100001010111111000110001011011010010110101111010111100010001010110001011111110000001011011100110011010101000000101100000110001001010100111011111100000000011101110011000000011110001111101111001111000000010001000100101101110011111010001110111110111111101101110001001110100011111110100001010011000000101110110110110000111001011001100110000010101110111011100001000111110100110001100001111100101110110010000011110101111100101101011011111111000001101100001101100001010011010101101000000000010011011000110100011010101001110100011100001101010111001110110111010110010100000100100001101000100000101001000010100010001011110100101110011011010000110011101010010001011010111000010101011100110111110111111000101101100101010110001001110001010010101111110010001110001111111010101101110001110111001100101101110111001111011000001000010100000101000111110000101010100010111010001010010001110000101011111000001010000001000010011100010001001000011110000110000011110101111;
assign EM[11] = 1024'b1101010100001111010100011101001110100101001010110100100010110111111101101110111000111101101110011101000010100010101000110000010101000100010001000100110000110100000011101101101110001110010110100010000100001000011010011101100110110110000001001100010100101111001000000110100111101000110101010100001011000110100110001101100011101111111101001101001111101011000100011101001101011000011110001111111110011010101010111100100101111011101101011001001010111010011110000001000000101111110110110111111010100111101000111110111000000101000111000011001100111101101001100010110001100011011000110101011011111111110010001111001010000111110100000001000011101011111100111101111000100000111101110111011110101011001001110110000000101011101011101011110010101001101000010000101100100000000010001001111110001110001011011100010010111000011010100000011110110000110111001101011010110111110000101101000001100010011100100011000110100000001101000010000111100101010100001111010001001000100011111101001010000010000111100101111001110001011100111111011010001111;
assign EM[12] = 1024'b0010011011111100101000100110101001101100111110001111110001100101110101001110000100000000000000001101010111001001011000100001111010001110100110010001101110000101100101011001101001111110010011110111100001000000001101010010101000111000110111011011100010000010110011000011110000100111111010100111101111001011100110110101010101111101000101100011001010110110000001110110111010110011111101001101000011010100001100110010100111001100010010011100111100111111010110000000101110100100110111100011110110010000101010111101101010001011011010011111010001001000110011001111011010000110001100100101101011011100000010000111010001001111010010001000011100001100001010111010110000010101001001110011111001010101101101000010100110001101111000111010011100001001011010000000100000110000001000010010001111110100011000110111100100111010110110101010111101101111111100110111010101010110000110010010101111011000100111000011010001001001000010111001101011111000110001101111010011010011111011101101100110101011010010101001010111000111000110010011001111110111;
assign EM[13] = 1024'b1000101010000010100111100011011001100010011011110111110001010110010010001101011000010111111110110100001110100011000000110110100111100110010000100101011101000101010100010110011001000110011010111001100111110011110001001101011101000110001111001011000001011100000010011010000101000100000110100111100111111110011100111110011110100100011010001011011101110100100011101111011100101010110101000001111011101000010000100100011011001000110100010110101110011000110000001010011110000000001100001011110000111000011011101100011101010101001010101101001000001001100010110011001001010101111111010000110110100111111101101110111101001000100101010110111000110100010011101110101010011100101100010011110100010100110010100010110111110101100100001110011000111101010100110001011111000000011000000001010111010000101000000000101101111110011110110011110110100001010001111101111110111101010001110111100000100011010111111011110110101111111000100000000111110111011001100100111000011001001010101011010001010101010110111011100111011001000010100101000000011111;
assign EM[14] = 1024'b0010011010110111011000110101101100000010100100100110001001010111111000100010011110100111111000010000100100000011111001101100111011001001000001111001001000111001000100001000101001001100101110000111100000001001000111110011110011101100101101000100011110001110100111101000000101111101101001110111010011111101100010101110001100010101101011001011001110000111011111011011101011100001100000000011001001111010100111010011110011101101100100111001010111100111001001000101001101010011010110000000101001000111011000101110001101101000100101000100100000100010111001100011110010110100111111011010001100010101001101101100010111001010011100111011101101000010000110101001001010000011100000100011011001100001100110110111100001010100100000100101000001000100111111100001111101100101101111101110001101110011001101000001100001110111010110011001111111100011111011100000001101100001011111100011101011010000101000101111111011001011101100110111101011011011100110010100100101110001100101011111101001001110011010011110100101001110101001110101000100110110;
assign EM[15] = 1024'b0000110011001001010011100100000101010100011011110111000110110110001101100001101110010011110100100101101011111000100111000010111100000110001101011101111010010000001001001111000010100101001011111101000011001011101100011000011011111001111011110000110111111100000100111011111000101001100010101000001100111011101010010000100010111101010000000001010101010110110110100111010100110010001101011001111010100110000111111110000101100011110110010111100001111111000010101010001110000111010000111010010100110101010000100100001110011101011110011001111101010100010101101011110010001100000011000000000001010101111111100001101110010001101011100000011001000011101010110001100000110101111100101101011110011000110110000010101111110001101000101010111110010000110111111111100110000000000000001011010001010010010010011111111101101111111011000011000100010001111110110000010100001111010000110000111101110110011111101110001001111101001110101101100101011010010010001010110100110000101111100110000001110011100010011111010011001011110101110000000111000111;
assign EM[16] = 1024'b0001000011111000001100111010100110110010101111010111010101011110010100010010111011001001010000011101000100011101011011110101110010110010101100111110010000011001101101000110001011000001110111100001000100111101101110111101000000111100010100110011010110001111110001000101010000110001001001011101101010001011111110000010101111000010011001011011101001010101011000000011010101011101110010011011101000100000110011011100101110011100110001110101000010110100101010111000110010010111100010000011111000010011100010100010110011010001110111100110101011011001010010111010010111111001100010011001110110110000000100110101011000110001111010010010011100001010100011010101011001110010100011011010011101110010001100001000100110001100100100011100011111010101001001110010110000000101011011111110110011111011110011110111111100110101011111010100011111010111110011011010010101001001011111101011011111001000111110110110001010100100111001000010001101100001000010010010001100110001111000010100000000101110011010101110110111000100000011100000111010111000;
assign EM[17] = 1024'b1000011101001101001010001101000001000111001011100111111110111000100000010010101101010101111000001010010011001100110010000101110111010010111100010010000110101101110101100101101100000100101111100101110101000000010100000110101000110111010010001011001101001101101000110110010000010100101101001100111111000101010111011111110110001000011111010011010011110001011010010000000000010000011010010010011101011000100110001111011101001000110010010111011011010110010111011111000100110010110101110101001000100111100111010101100000000100110000111001100100010010111011101011101100000011101111001111101101001010100111000101111001010100000011110001011110111000101000010100110011100000011110101000001111100011101110110100011000100001111001100111100111100010000011100111100000010001000110110111011010110011101110101111000100101001010101110110011111110100110001100101010000111010010011110101001011111100011011010010111011000000100001111110111001001100011011011110111001110110010100111100110011101111001001010010011100101101110000100110110000110110;
assign EM[18] = 1024'b1000010001011111101000101101101000001100111010111101011011111000100101100010110101101000101100011010101000001000100110011010010100010001011110100100100110000101101011010101001011101101100011111001111101101000000000000001010101000101101101101110101111101101101010110101011111110111110110001000101010110111101011011101010010100110010010011010000000011000101100001100010001001101000100110110010101111000100111111111110111010100100000101101000010111011110011110111000110100001000111111110001111000001101110000010000001110010110001000100101011110101100001110110011001010011111111000110101001001101000010001010000000101000011100001000110011011010000011110001000001100110010101000101011100110010101000100111111110000000011010101111101100111101001010100100111100100010111011111001010100111001001101111010000001011101011011011011100100110111111110010000000001110001010011000011110010101111111000001111001001010000010110001011101010011111001000011110011000011000011001111010011110101010010111010001010111110111110001110101001000111111;
assign EM[19] = 1024'b1000011110011110110011011100100110001000111100011101010001110111110011001100101001111001101010001001001010001010111011101111001000011000100000011100110001101100111110011101010110010011011100000000101010101110110001111111101101111010111001001001101110100000110000101010001100001101000011101001001000010001111111111010110000001110000100110111011101110101010001011100100010001000111000101010111001001001110000110100111010100000111001000111001011000111001101111101111101010111010011011001000110101100001010101101000001110000011011110001001110011011100011011111011111110011111010001110100110000100111000010100101000011111011100000010011010101100110011001000111110100011000001100101000100000001110100011010010100000110100110000001101101100101101100010010000011101100001001110101111010010101001010000100010110111011111100111001100101101011010010111011111010011110011101111000010111110100000011110111100111111000000100111001001101101010000110101001000110111001001111101100010101100100110001101001011010111000110010100010010010100101;
assign EM[20] = 1024'b0101100100111100010011001001001001000001001010100100110010000101010111101010110110101100010001110100011111100001001111010111001111010000001001000000010111011110110100011010000110101110100111011111010010101110101001011001010010011011011111110010001101101111101010111101110110001001100110110000010000011010110001111100101001011010010101011010111100111100110010110010011111101111001111101110001100111100101101001011011001110100110100001011111110000111100010110000001011101010000010111011001100010100011011111111100001000010001101001111001000011000110010100110001000101101001110101100100011001110111100001011101100111001010101001100101101101001000110000110100011101011000011111000100001101001101010011010011111001011011010100100011111111011100000101011110001000001101100001011100110011001101111010100000010010001000111001010010101101010100001111100000101101000011100000001001110100111000110101011110111101001001011010010111010010011011001101110001101100100000010000101001110100011110111011101001000100000111000101101101101011000;
assign EM[21] = 1024'b0100111111100011111111110010010111001010111100101000000000111010100111000110100001100010000111000010100010111000011111111111001011101101111100110010111110111110110110010001111100110100011101000010111010110101100100111111001100101111011001001110011100010110000000000110110011111101111010010111001111101010011100100000100111001101001000110111011011100111000001110000111110100001011001011111101110011010110010001000101000110110001111101101001111111110000100100101100110000010101010111000000010001011011001111110100001100111101010000001000000101110111100000001001011011101110001101110100011110100100011000000100011101100011011010101011100111000000000100000011010101100110000111010001100111101000101000100010101101100001100110110110010000011110111101111000110001101101110101001100000000001110011010110010010111101100110100101111110101001110010111011001100011110010100001110100001111001010001001010010000101100011100010001110100111011010000101010001100101000101010100101010110111000000100100010011011010111010101100100110000101101;
assign EM[22] = 1024'b0110011011111000100000000001010011011101001101010011111001110001001000101001101110001101010111110111010001010101011100001100101111010100000011011011011110001010011011100111001101100110011001001011110100101110101011100100101001010001111101110001010100010100000010101001000001010110010010111111111000100101000000010111011111110101110011111111101111000100000010001000101100010001010001111110011011010100100111110100011000010110010011101000010010101001001100110010111111110101010010010100001001110010101000110010011001110101111100100101100110001110100100000000111110000111000100111011101010110100010111000001101100010100100101110100100011101010010010111010000001101111011001011000011101011101100111000010110111111011101101001011011001100010000000001011110011100011010000011001011010011111110111101000101011000100111011000110101000110111001010001111010000001000101011000010110011000111001010011011100111011110010100101011000001100000001110011110011110010110101000101001101101101101110111110100000010110101101011001101111011100100;
assign EM[23] = 1024'b1100011111011111111100111110101010001100010100010001011000100011111000111001101100001000001100111110000110010010111001100111000100101000011110011001111111010010011000111010001110001000010100000010111011001001111000100010101111001111010010010000111010101101010000100011111100101100110100100100011000100101001001001101110111011101110110101111011101001000000011010101100110101100111010100010011001110011101111000110010000011111110011100101000110001101101100100000110110000110001000010000011110100111001101010111110100101111000001000101001110001101010101110100001101100100011001101110101100100001100011011100011101110111100111100011011111010011011010111110111010111000010011010000110010010001001100111101101101011110010110000011001000000000110010011011000001101010110111011001101000111000111011111001100100100100100000100101101101110010110000010000111000101001110101001111010000000000111101101101110111101000000000100111011110110110110100010111010100000001110111111011100001110110110011111111100111000110000101010000101101000001;
assign EM[24] = 1024'b1011100110010010110111011010011011011110100110110100001111100110101010110110010011000011001110101001101111111000000110000100011100011001011000000110001101100000010111101011001100001000100100101100010000111000111101100010111101011000000000000010001011010100101111111000111101111011111101111010001001000110110010001011001101100001011101011110000000000110100111100000110000001000101001100010010011010010111000100110101110000011100011111111100101110101110000101111011000011100010011010010100100011001000110100111010101010100101001111011100111000110110001010110101011010100101010101010000000101110101001001100111110001001000001000010000010110011111000000110111010110111111011111001101010011001000101110111101110100110011110010100110101100011111101100011000101110001001110011100100110110011110001011011000000101111000000001111111011110111100111111000011110100011010100001010100010010110010111011010010011111111010010001100100101111100000000010101001010101010010011000011101111001110111011001010011010100001011111101000001010111111;
assign EM[25] = 1024'b1010001101100011000000001100000111000111111110011111011100011011010100100111001111011101010110010000010011100000000110001110110101011011011000110010111110010100111110101001101101000111110001001110000000011110100101001010111011011111010101111001110101110101101110110001000010110011101100111100010001100100100011000000110000100110010101011010011100001110100101000111000100110110100110111100011011111011010100011101101001100101011110111010111110100011000001001000001100010111000010010110100000011000000101001010101010100000000100111010111110011111000101001110111001011000111101000011110100001101111101100111000101001000101010111010101000000111101000110011010101110001000101001011101001101001000111100000101011000110011101011000010011101101010001001010101110111010110011011000011010001001101101011001010110001011111101111110100000101000101100001010110101011110100010010001011001001001001110001110001101111000000101001001011110010100101111010100000011111011010110110111010011111011010011111000001000100111011000100011011011101011;
assign EM[26] = 1024'b1110110000100000110110010100001110100011110101100110011110011100111000001101010001000110010101011111011101011100011101100011011101110110101000100110101110010011001110101011101010111001100100011001101111000001111111101101100101111110011000000001010111110110111010010001110010001100010100110000111001000000111010110000100010111010001101110010001100000111100110010000000101101000110101111000001110111000000101001011001111110010011000001110101101111010100010001111000000110000101000110001111100110101001101001110110000110001111101111100110011100101111001111100011111110011011110100111000110101111100111010010011100001010110001001000001001111100111001001101011011110000000100101010000001100111101101100011100100101011001101101001101101011000110011000011100001100001100001101001101101011010011100010010100000010001010011101010100100010001101111010101001011111010111100010011010100110101111100000000111001111000100110111110001011001011001001000000010110011110101011100110001000010111101101111000101000010100101001011010111100001110;
assign EM[27] = 1024'b1000001011010010111000011111011111100001111100111001011000001100110000000101111100001001000001101001010110101011010011100001100001111001001101000100100010111101100010011000010111001001000111001011110011101001101001010110100111000110011011010011101000101001101011101111010001001001100111010100010111111001100011100101100110010011111010000011101011111111100111111110001101101111001010101110001111011010101100100101111000000101111001101000101001011111001000000110000101001011110010100001010100101001000010110111100110110110000011010000100101100000111001111100111010011110010101101101010100100101100100001001100000111011101001100001110000111100001101001000000010011011110101011100110011001100011011000110110000001011111010010011110010101011010011000000101100100001110100101010100000111101101001011100111000100100111010010011100011100101011110100001101000101000100001111011000010111011010011001010010011101111010000000100101111011000110111110101111001000011110110101011011000110000011101111001001011011011011011010111100010110011;
assign EM[28] = 1024'b1101110101011001011000010101110100100001101011100100000011001001111111111111101110110001011000101001100001011110000101101100111110111001110001101110010110010111110111000010111011001111001100111000000110010000100010111110010100011011101000000000101110101101010001000001100111011111100100110110000000110101100001101010011111001101011000111001000111100101010100010000101111011001000010110111101001011000110010011011011011010100101100110001000100001001111101010011110100001011000100100001101110011011000110110011001110001000110001101111001010001101000011110111100111010000100101110001000111010111010101111100001010000111111000011100100010101110111100110101101011101001010110100111101011010110100100000001000001000111100010001110111110001100010001101101110001110100000010100111001000011111111111100111010000001001010100110110101100000101101000101111101000010011011111101011010000000100010111111110111100101110001011101111011101100011011001100111010000010011001001011011010100000000010010101001100001001111001100000101110000001111;
assign EM[29] = 1024'b0010101100011000000001100111100001001110110000100110100000101011011010000110010000000100100001100101111010101110111000001100101010110011000110100100011111011111000001100111101111001101100001100000101011110111111101001110000110001110010001111110110001001000110110011000111010001110001100000000101011001000011010111000010010111011000000010011011110011010000101101000010101000101111011101110001000111010011011111111111011100000011000111100101010001001110111111011001101111000111110001111110111000100101010111101010001001110001100110110110011110101111001110001011110001110110000100001100101010010010100001010111011010101010111000100101110011111110011111000010101101100001001100110101110101000001100100101010000111010111110100000111011010110000110111101100000010100101110001101001001001111011000000010100110101000100111101001101000100101101011101010100100011011010001111111110110111110100111000001100001001100101100100110010000101011000110010101101010011101110011110100011100100010001011011101001110011010100101110010011011101100;
assign EM[30] = 1024'b1011111000111101111001001010010101101111110011011000010011000010001110111110001010010011010011110100101011001010011000100111011000000111000110011001101001010001011111000110010111000111000000000000001101111010000010101011100000010111110110000001011111010001110101111010000111110101101101101100101101101010111101001010011010100111010001100000101101001011011010011101010101010111000010000111101110111110011100000001001011111010110101101110000001111111101100000000001101111001001001001011111010000010110111110110111110010000110111011010011100011101101011101001100011001100011100110001101001111011100001000010000000010110101000010110110000101010110011101011010111101001010011000001100110100000010000001110111000011010110011111011000110001011110110100011000101010010001111111110000111011011111000111011111110100100011000010000010000010011100000000000000110000001000000001111110011010111111101000111100010100110111101011011111100001000010110111110111010110101000001000110000000010000101001101111001111100100001111101101101001111111;
assign EM[31] = 1024'b1001101011101100000001011000100001010000101111110101011100100010101101100010100001001010010010011101111000110101000111000111010000001101001110010001110110010111000110011010001001101010110001000000010110011111110010011111101000011101111101001110000000111100100011000110100001011000101011000111101011101001001110001001111100101111001000100101010100101101010101010111111110011100101010011001101110001101001111100100100011110011110010111001000000111101110111101100001010110001001111110010100110001010010001111110111000010101111101111001000100001111101100010010001101011111111111100100100100001110010001110101001110101000001101011011100111011100101011100010010000001011100010001001010001000101010100110100111000001010111011101111011100100100100110101100111011101001100110010111110001101000001110011100110101011100001001110100011011110011001111110000101111100111111110101001111100110000001001010100100100111111000110000100000100001110000101101000100010110000110010110000001111101110010111000010110011111010110100001001100110100001;
assign EM[32] = 1024'b1101010100111101110111010001010011111001011010111110101110011101000011010011101101100011100101000100010010101000110011101010001111000000011000110110110111100111100001000100001010011111001011110110000000001010111111011011011110010010111100000110010011101110111101101001001000101001101011001111010111111100000100010110000101001111011111100110111010001111011000000111010110010111101011000111000000010100000000100010101110110001101110110011101011101111100110000000001101101010110100100110010111100011011001010101011000111001110100000001101111000010011001001110101101101000011001000101011011101101110010101111001000101010110110101011001111000001100110001110000101000101001011000011000100110101011110100101000110111010011010011101011000110000001010110011101001000001001111011111000110110010010000011101011111101110111111101010111011110011010000010111000110110100101010001010111001010101010110100101000001110010010010011100010110010110001010000101010100111011110001010000110001001101110101010000100000111001001000110000000101011110;
assign EM[33] = 1024'b1111111100101111001001010011011101101100100111000100011110010000010111010001110100101110110010011100100111011111100000100000011011100010011100100000100100101001110110110010111001100100000100101111010001101100110000100001100111000110000011010111100010001011100100001011010111000111101001010111110110110001100101101101010101000011101001100001111101110011001011011100111101000111011011010110110101100000011000100001011100010101001101011101101011001110010010000110111011000100001000111110000110000100111001000000010101100100110101000111000001101110011001101010000101000000111110111001001101011010111000011100001000100110011001001100011100011001001010101000110001110111111111000110010101101110010011110101100101100110111110000110010010101011100111100000010011010111001000111101110001110011000100001111110101101011111000101110110001100010111110111000101111110011010010011010101111010110100011000101010011101001110110010110111101111010000001100100101111001001000000101100010001011001000110110011100010101110100100110111010001001001;
assign EM[34] = 1024'b0010001011011111001000011011010100011011111010111100001010010110011101111001000110100111001101010001001101011010100101000011100000111011111010001000001010000101010110001111101110001100111011111110100010100100000000011011101011100000001001101010011100000100001110101110011100010010101100100110101010100100011110011001110100110100010000000011010010011010111101000111010111010001010110000011100000101110011000110011010101000011101001011110110010000000010000100111000001010000100101101001111100100000000101111111100111011011011100110111111001100111110101010101001110110111100101110111100001011010101100010010110101000111001011100000111110010011110101010001110110001000110110111001110001001001001010110011011100101011111101001010001111110011010101001101111101111010101111100100100110100010101000111100100010101111101111111001000101000110000000000001011010001100110010100100101111111001010101101110110011010010000111001011100001010000101000110001110111010101101100110110000111001001100100111011000100011101000011011111011110010011;
assign EM[35] = 1024'b0101101100011110010000111100000110111110111011000011000010000100010010101010100011100010010101010001010001111000110110001100111000010000001000101000111110000100000100001101111010010001100111001010001110001010001010110100101010011110101100010100010001110001100111111101011111111101010100111101011010100101110101000010000001001000100100011110111001100011011000000111001100111101011101110111010111011110010001100011110010100111000111101010110110000110001101110000101101010101001111011001101100101000100001100100101111111100011101011101000110110001101010010011110100011100110010011111110001110010100101100010111111001011100101010111110110010010100010000101100101110001111111110011110000110111011110011000101110110100110011100101000101010000111101000010011010101111111111110001000101111111100010010100000010000110100101110001010011011110100010100111110000000110111100010001010100101011010010011000001100100111110111110111100010010000000001001100001001000011111101110100101001000100011100101100111101111010010100011110010101101001;
assign EM[36] = 1024'b0100010110100000011110001010110010111101010100000110110110011101111110010011000111101010010100100111011001011001001010100111000011011100010111011100100011001111101010101011000011100001101101100110010011001101000011111010110010000011110000100111100110001011010001101110001100111111011101010001010001101110000100111100011111000110110011011111100001101001010110010111100000101111111000100011011110101000100110011000010110100100111110100010111101000110100110110111111000011111001110101111001011000011010011110000001110111011010000100100101111100001000011110000001011110001010101000101001000100001001100011000001110011101100110001000010010111001111011011001011000011010101000011100111000001000001001111011100100111011100000110011000011001101000110100100111110001100001101101110101010010110001110100001101111011100011101101100110101110110110000101010000100010000001011101010001100111010001110011001010110111001100100011011111100100101111000010100111101110111001010011101010100011000001110111000110010010100010111011010100010011001;
assign EM[37] = 1024'b1101100000101100100101000110001111011011100111000101101001011001000101100010001100110000100011000010010111011111100111100111010001111110010110001110000011100010111100001011100001100111000110101001010101011101111011010000010101011011011001100010100001101001101000010001110110110110101111010101101000100111101000011000110000001011100111100011101101111101011011110011100101101010110100000010100010000011101100110010100011100011001001100111101001000110101011111111001001100001110100110011001110110100101001000010010101010101101101111011110010011111110101111101010000001110001011011111111100101000011001111001010001000010000111010100000111100011011110100110100000011100010111111010001100110101111011000011000111101101010010100100101101010110100101110011011011101011000111001001010100000010111110001110010001001010101011110011001010100101001001001101011011110111000011001101101001000001110010010101010011000110000010101101011100101111011001011100000011000010111100100011000100111011100100011000010010111101010100000001101011110001;
assign EM[38] = 1024'b0011111110111001011100101100010010011010101111101111000100001010001101011000000000010111011001101000111101111010010100110011001100100010101111010110000101000111000001000110110101111110100101110101111011001011101000000000000010010010010011001111001010011010011101011100100001011011101000000110110011101001011100011011000000011101011111110000001100001010001011010001011100010001101100000001001010110111100111011110001111111101110010111010101010101000101001110010110011010101111111110010110110011011101010100110011110001111111100010010011000101100101001001111101111110000000000101110110010001001100010001010111001101111010101011111100010111000011101000000111000010111010001000110010011101011001110001111010101101111010100001111000111101001111010000100001111011101111011111111110110110100111000011100100010001010000101101011111010001000110110110010110001000100001011110010011101100011000000001010000110011101111011011010001001001110001100110000100101111110110101000011011001100000000110010100100001100100010100101010101000110110;
assign EM[39] = 1024'b0111101111110001100011011100101000010010000110001001011011100101100101101011010101001111010110000001110101011010011001010110100000001001001111110000000100100011001010110000010010100010101100100001111101101110001111111110111101011010011001000101110001000111110001100110000100110010110101111110001110111110011001011100101011010110001101011110011000001100011110010001110111101011101000110110101010001100001100010010000011111001101100100010101001000101101011101110000001010010000000101100111101011111001111101010001001101100000001001110110110110110000011100110001010100011000010100111010011010110101001101000111100010100001001100111010011101001001111010101110100111100110111110001001011110011001010000110000001010100001011011100001100100111110011010110110101010100101011100100111111100100110000111010111011010110111110110110011100100011111010111100100001001011001101011111011010111000011100001011010000000100011001100110010100001001001111111110110001000001101111001000110110100100001100011000110110001110000110010010101011101101;
assign EM[40] = 1024'b1001100100111000111010001111100010110100110101110100010100001001111110010011101011011000111010101101110011110111101110110110100011000010101001010011011111110010000011000111100100100011010011001011111001011100100011111110000111000111101111001100001101010011011100101101000000011101110110111111010000110101111101100100111111001111100000001101011010001000000001110000100100101101100010100100000100000000111000100011111110101011111100101111100010011100110101100010001011001010011010011100000110110011101010100101111100011001000110001110100000010001101101110110111000110000111011011011011000111011111101100101110100101000100000101111010010011101000110110110111110100001110001001101010101010011011001001101101001101111010111010000100011101110010011010011110001001000111010010010010111111000001111100110011100110010010010001010010010101001000000101100110111110010001101111011100000000010010110101101111100110000010010010010111100011110000011110000000001000110100001000101010100101010100110101110100010010001101001110100101101100101;
assign EM[41] = 1024'b1100000101011110100110000100101000100111100111000110111000000000110110100001111011111101101001011010100010001100001001001000010011111110110011011111011100011010000110101110010011111100010110111000110101001010010111010000110101101000011110111001000011011010000011111011011001011110001010101000100100000100011110011101110101011110101111100100010011001001101101100001110011110001111101111100000111011100101111010010010000010011011001001000110111010100010110111100101011011000100111000110011100011001100000010011111000110001101001011010001011011110011110000010100010100011101000100101010100111000010010001001110100010011101100011110100010010111100001110111000110011110001001111101010110101111110001001010000100000010001100000100100001000110111000101011111011100000010111101111101111010111111100011010100100000001101101011000100111000011010101011111000010111101101001001110111110011111111001110110111010111001101110111100010110010100100110101100000001100001100010000111100100011110001000100101001000010110110111000110101100110000;
assign EM[42] = 1024'b1001010100100010101011110000001000011000110110001011101101010010001110111001001010111110000010000001010110010111100101100101001000001101011101100110000001100011110111100000010001010110111010110010011101101010000011111001011000111010100000011011110110010011111000011001101110011111000100100101010001010100011100100010011111011010001011100111110111011100010101110100011100010001010011101100111101001011000101101011010101110100011001111110101101101100110111101101011001111011000000011010001010111111101100000101000000111010100110001011110000100101101101011101010010100101100101000111111001011010010000001010101100101111011011011101011000111011001000011100000110101001101011010101110111111101111011101110111111110000100010011011000010100001110000100110001010111000011000001001101010101110110010001111111110101110001100001101100011001101100101100101011010011101110101111110100111101101010100011000010010000000010000110010000101110001100000100111110000000100011001010000001010111011011001111111110000010101100010100111000110100100;
assign EM[43] = 1024'b0101011100000100101001111110010000000001011101000110011001010101011111000000001100110110101100100111011001011001100010110001110011001110001100000011000000011011111001111110000011010110100001001101101001000110010001101110010001100101111101101110101110100000001110110011111111011110001000001101010110110101001000111011001011101101111000101101101010100000000111000101001111110001101010001000111000010110111110110110010110000111101001110111011000010000101110111111101001111110111001011011001010000110000011111111001010011110011110001100011000101010000101111011010100001011101111000100011011101000010111000000011100100010010000111110011101110100000000110111010000110100011010111100011111000110001101101101101001111001100010000000110101001001100100110010100100101100110100101011111000110111001010000010000001001000100100000100100101011011010110011001110011010010101111000100001110111000011100001101011110110001110001101010011110010101110001111011011100100111011000110000111001010011000010100111101111110100111001011111100111111000;
assign EM[44] = 1024'b0110010101011110011111010100111101001101000111001001101100001111010000110100111110101111110110011100001001100011110101100010000111010001011110111001100000000000000001011101101001011110101111011000110001010000001100000000011101110111001011010101011001100100001000100110101110011100010100001111010011100101111001100001100010010000000000100010110001001000011101010111111000100100110101011111100001101111001010011000000011110011100100000100010111101111111011101001101011010001101100001111101101101110001111010110111111101110001011010011110101111010110001100010100001111011100011100110010111001010000110010101111011111000011111110010011001100001111001010110010011100000110110110000111111001110000111001011011111011000011010110101010111010100000011101001011100011011001100001101101000100001001001011010100111001000000000011110111101010111010000000100001100101101010011110000111111100001111000110001000110100111101010000000100001011001010000110011111110101111111000111111010010110100100001001100101101000110001100111100100001000011;
assign EM[45] = 1024'b1110100001111101011101101110011001101101000111001100110111001011100100110000001011001000110101101100110010000001101110000100011110001010001001001101101011011001011011100000101000101011101000110000001000001000111100101011110001100010101000111111110110100000100110011000100001111010101101001001111111000110110100001111010110001101011010000110110000010001101011100101010110100101010010000000101001010110110111011001011101001110101110000011000000101001011011001010111100000000110000110011100010111011010100110101001101111111010100111110010101100110100101010000110000011011011010101111101110101000011000000110011100101110011110111111011111001101001000010101101110010000100001000111101110010011100100010101001110000110110000001100011011110010000101011001101111110111110011000001111100100100010010000011001100110111100010101010101001000111000111110001100001111111011110011010101001000111000011110001000110110101100101110110000111111010100100101111011110000111001110000001111101110100111111100110010101000101010010110010110100010101;
assign EM[46] = 1024'b0001110110100010011011001011101011010001000010100011011110110001100111101101101100101011010011011001110001101010110010000100111101110101100010000111010001000111010111111110101100010001100000001001000010001010010010011100010111010100000001111011100110000000000101101011111101011001110010101110110010101010000101010001000111010010111001101100010011000101111000001000100001101110000010000011100100010110111101101011111001000101100011111101011011100000101000101111101101011101011001001101110010111011000001011000010111111011111001110001011010010001100110000000111000011111101101110000001111000110001001000000011010101110011110101000010110111100111010000101110001110011011110000001011010000101110000011101111101011111111010110011000011001101001011011000111101111111010110011110101101101101100101101001110111010001110100010010010010100110000011001011010110001011100001010000100101101110011110100001011000001010110000110010000000101101011100101100011011101100110101001101000111111101111011111011101010011010010000101011010010101000;
assign EM[47] = 1024'b0010101100111100000100110110000011100011101011111101111001110111100110010101111000110000110010101010101101000111111100100001110101100000001110110100000011001110100110001100101100001101110000100111100000101001001000000000010101010011010000010101101101000011011110100001001011111101100001111111001011110001101110110001100110111110000110001000110110000110011101001101010110101100111001111010001111100011010010000110100001100110011010010110011001011101110110010111111110100101000101010011000000100100100010111001000111101110111101011101101101100100111111101011000000111110011101110110100010110001111010111000000011100101100010111011011101000100000000100000110101011010001010010110010001010001000001110100001011010000000101100011000011110101011111011001001110100100101110100001101011110011110011011010110010100011101101010111101111011100000111111000011000010011000111001110000001101001100011111101000011100110100100110111010110000110101001010011111001111100100101101100010001111010100000101100101111110101001010001000100111011100;
assign EM[48] = 1024'b1011000111111001000110111010000101100100010010011111010010000111110001000101001110000000110011001100000001110101101001110100001100110000001011010000011101000001101100101000010111000001000101100110110010101011111111000101110111000010101001100000000110110000100111010111100100100100100011101101111011100000010101100110000001100111001010000110110100000110101100011010011000011101011110001010110100001101101101010011110001001111110001110011000010001100111110111011011110010000001110101001010111101111001001011111001001011000101110111000001011000010110101101101010001010001010010110110011000111011011001011001001000000111100011101111001100101101100100101001101010101010111000001010101010101010111001000100010001001111001110000110111110011100110001110110010111100000100010111110100100111100111011001110100000110110001110100111111011101100110100101001000110001001011110011100110111111001110001101101111001110011001010011101011011110111110011100010100000111111111100100011100111110001100000111101011010000111001010011000011001011001;
assign EM[49] = 1024'b1011101110011110000001011111110010110111011101100100001110101110001010111110111110011101011110011011001100000000011111010011000011010110011110110111110100000101011000010010000100001010001101001011110110111011011111111000011011000000010101110110110100101011111101000110111110100011010101100001001101111110100111101110110011101001101011101010011101110011000101001000000000010101001111001100011010111101010000001011100101100111111000101000011010011100001011100101010000100100111101000111101010101001000000011001100100010110111100000000111010010101000110010101000001000110110000010110111001111011010111110110011101001111011101000100001001000101010011101101111111100000010010111101001100011101011011000110000000011110100010110100001101001111000101110111000011000011101011011000000011101010101101100100101001110011101100010000001011011010011000011000000111100001000001111001010001011000100111111101001110011001001001111011110101110011010010000110001000001100111001001011011110111010000010001000111010000110110000111001110110000110;
assign EM[50] = 1024'b1101110100101001101110001011100011100011110111100111101011001101100010110001100100010110011010010001001011110110001110111100011111001110000000101011111001111110100010011100011001100001001000011100111011010100000101101001001110011111011001000001100010101110010101111000111100110001001001101011010110100100111101100010011100111101110100110000001010110111001011001111010100100101000001100110111110000110010010111010011001010010000000110100111010011110101010100010101010001011001111100110110111010010110111000100000110011100111010110001001111010100000000110000100111110111111101010011001000011000111110011011100001100100011101101011110110001001111001001010010001000000010001001110000010001100001101100100101100100101001101100010001111000011000101010101011010101100111001010010011111111100111000110011111110001100001111110110101110010101001001001111010010010110000001000010101011000110010111111110101110111010000111001111011111000110011110000101110000101000110111110101110001111000001010001001000011101001111000100010010010110000;
assign EM[51] = 1024'b0101111110101100101000010111100011100010111001001001111111010010100010001001001001100010001010011010111010011001111111010000101100110100010111010101010110110010111100000110011110100111001100101101100111010101001110110011001110110100101100010011001111110011101110111111000010000110101111011000000001000101110110100110001011011000000011101001000010110001010100010100000000101001110110101111101101010011010111011100011000001011001100101001101000010010100101100001011010100100110000110110001110011101110100111011010111000100010110110010001100110010100101100010111110011110100000110000110011010101101001000100100110010111010110111000000011100001110100001000000000111000000111100100001001100110100010101101110100011111101110110011000111000111111100110000110000001000101011100100001001111111011110111011100111100011110111111110100111110011011111011000001111110000011110010110100011110111110000001010110101011100111101011000101100111010111100110001001011110000001010100001110010101000100001010100001101100011100001100001010101101110;
assign EM[52] = 1024'b0010001101110110111101010000111011110100110010001110111110110111001010001011010001001001001001110010000010100010011001000101000010100001110011000010101101010101010100000011010111110110111010011101100100000010110000100101000010011100010101100110101010000100111010111000011101100111001001010110100110000011011101010101110110110100111011011111011101100001101111011010110001110100110000011100000101001101001101101010010000110010001100011011000010011110101001111100110110111100000011001011100111010111110011001010101010101001010001010011111100011010000000011000010000000101111100110101001111000111011111010100011100000110010101010010100011011111100110101100100101000100100111100000111111100011101001111100110110001011011101100100110011001111101100010010101001100010111000001110111110110000101010011001001010010111001000101010001011100001110001110111100010001101110011110010100100100011100100110011011101111111100101011110010010011011011001001100101010001011111101011100101100010010100011101010110101110110101100101000010001010110;
assign EM[53] = 1024'b1110100000100010011111110001101111001100101110000101011110110111011111010101001101001000011000011100001001000110011101110000011111001101111100111011110111111010011101101101000010111111110000111101100011011011011100000000110000110110110010010010111100100011011110111101100101100100101111001101110110101110010100000110000000010001111110110001101000001100101000011000001011101110010100111100011011010101001001011010101001110110010101001100001110011101011001011100110011101010010010010110011011001011010110110000111011100100010100100000001101001110100010111000110011111100100111000110101101111100101000110010110010111100101011100101110111011111111100111011101001101010001011001101110101000010000000100111001011101001110010000111010010001000001011111101011000100011110101011000110000001010101100011000010000110010000100010010101000101101011101001011001110111010010110000101000111110110111010100011100010110000001000010111010001001100000010100001010101000001110000110100010101010100101000100100001101011111111110100011000100110111;
assign EM[54] = 1024'b1010011011000110100000010101001101101100111000000110010001101110101010001010011011010111110101000000010111010010110010101100000110110100011010010000010111110100011100100010111111010101011111100000001011110000100011011110101111010101001000000001111111111100000101010100101000010111011011110000000001000111001110111101100010011101001001110001111111000110011101000010001101100010011001110000011001000100000101000000010110100010000010010101010101010100111111111010101110010011101010001101111001100011100101111010110011101010101001010100011000111100110101111000011100111110000111111001101110110001010111111011000111111100100000101110110111101101000001100010111011100111000011101001101010100011000101110110111010001010000010011100010010101000111111010001101111101101101011011100000111111100000101010000111011011101101111110110110000110001100000110011111101011001101001000001101110111110001011001011000101000101000110001100100001011011100001000011000110111011111100010101100010000100100110001111011110010000001000000111111110100001;
assign EM[55] = 1024'b1110001101000001001101110100110010110111001101100011110010001101101011000111001100111110110111101111101000010110010110001010010110111101011110101000101100010011000001010111100000110010100101001011111111001111110000010011111101101010110001110111000100100111100110011000100010101101010101001001111100111000000001101001110101000001011110000101110001110011101110111101010010000010110000010011010000110001111011001100111001010011110000000101111100000111111001000011110101010111101101111110111110111101001011100001011000110101001011000110101110001010010110110101110101010011110110011110110001000001001100110001011100101000110111111111111001100000001111010001010000110010001001110001000011001000111011001101100010100101111110101010100011110111100010010010010001100110100000011011011111011000010100100000000101011110000110010111000000011011000011110100011010110100010110011110111000010000101000010001111111110100111110111001011000100100110101000110010000010011110010010001100001000101010000001101011110011001110101011010010100100001;
assign EM[56] = 1024'b0010110111000000010101011100011100000011100011100111100111011010010111000111001111110111100101111110011011100100000001101100000010000101101111110110011111101101011101111101000101110100011010100000110100000010111001100011110011100111010100011101111111100111101011010001100110011100001010001110100111001110001000011010000101111010100001100110001011100100111110100110100101001100101010000111010100111101010101000000011010000001010011010011101011010011011100000000001101010000111111001100010111000111110001100010100100010010010010101000010001100010100111001001100011111110011101010000000000001111010010110001100000111100010101110100100110000110111011111001010010111000101111011111011100101100101110010111010111100000001111001001010000100011000101100011011110011011101001111010100010000011000001111100001111000110000101101000110000101110001011110010000100010111010001010100001011011010100001011111101111000000010011110011101100111110110101101110111110011101011011111100000110011001110010001000101100110000000111111100011101111100;
assign EM[57] = 1024'b0011110001110001001010011101101000100100110111100001011000101101100111100100111000100010010100101000100111100110111010111000111010101010011110110011001001000000100000000101010101011001101001001100100010101101110010000010110100110100001011010110010101010101001010011000001111111011100110011010110000011000101001100000010100000001110011001110101000010000011110010110111000110111000100111001010100101110110010101001111111000110101001111100110110110111110000111010110100111011100110100010100011000000101101101010001111010111001011111000011011010010001011101100101000100011010101011110100101101111111011011110011110101101000101101000010110010100001110111000110110100101111100111101010100001101010001000000011011011111011101000000001000010110100011001110001011011000101110001110000001101000111100111111100100010110001110001111100001110100100011111001111110101100101100110110110110011100111100001110000110010100101111111110111110010100010100011001100110100000110000000001110000010111110100111111110010011001100001101101000111100011;
assign EM[58] = 1024'b0011011110111101001101111011001001111010101001010111001000001011110101001101111110001100100110011100110000111000001110010010000100110100001101010100110110111001110110101010110000111100111111100101101101001001000111000111011011001001000101101010110111010111111001001101001101000111000101010001110110000110100000011111100101000000010000110010100110001110000011011001011000000110111110100111000010001000101111110100100111001010111011000111000111111011110110011101110011100010000011000010001000101110010101011110011011011011000111011011011001001100110000111110111011110011001001100111010001010110111001110010111101001000011001100010111111101100000001111001011111000110011100101011101001010110101100001101000010011100001011000000000010101001111011000101111001010100000110101000100110100001100011110011011100010101101100011100010101111000001111010011001010001100000001000000111001000111100000111011101100010100010100010111100011110010100000100001100111111100010100101100101011000010101001111110111011001110110011100110010101000110;
assign EM[59] = 1024'b0101010010011001110011110001010000011111101010011000011001110010010101100111011111001001001111000011001101000100110011110110001000100111111001111000110001000011100010110010010101101100111101100100110111101110010011001001001001011100110111110000111010110100111010001110000010010010100010001111110000000010010010111010100010110100001001101010100111011010110110010010111101111101111100000100110011101010101110100110101100011011111001010110000110010001101100101111110100000010001010101011101000110100001110011100000111100111110000000100110110110001111011010011111011101111111011010100000010101111001101000011100110111100110101100011010000010110001011001101010001010101000011010001011010110010111011011101110100110000011000110101000001001100111011010111010001011110011101100000011000010000110001111001001011010111100100100001111000001101000000101010001011110010101100100110001111000011000110010001101001001001100101101110101001000001110111101110101101110000001101110010011000101011010111100110010001011110010101100111000010111111;
assign EM[60] = 1024'b0101001110110011111001001011110000111011111000010110011001011010111010001010111001001011111101111010111101011111010100100001100101011001110100011000010011010101110111001010111010110110101101001100000100001101111010110000010110001001000111100100000000111011011101001100011111011001000110000100100111010010111110000010111010011010000100111000011000110111010010111011111000100100001100110111110001100000111111101011000101111000100101001110101111001010101000010001011011110101001111101101101001111111001000101100111011100011001011111010100011110000000111011110000011100010100000001010100111000010000000000111110000101000010010010100001100011100000001001001000010100111011001111001110010011010011111000100110010111110010011000111000001011111111100010011001101100110001100011100000001000010101110111011111101000111100111001010011001100101101101001011110100000010111010000011111101110011100010100011001001100001101101110001011111101001111001010101001010110110001100000011111100101010100111000100000110010110110101100110001111010000;
assign EM[61] = 1024'b1101000100101010011110100011100011001100110010000111111110010100110100110111100000101111001010000101101011001011010010100110101110011000001011111001101010011100011001110000110001101100011111011000111101100110111000110110101101101010010100100111110001011000101010100001000101111101001010010101001100001000011011000000101110001011111011000100110101111100000001100001000011011101110110001110111100011001101011101000110000011011100001111001000110000001111010001110011001011010101110000011010010010110000110010011010011100101011101001000011011001011011011000011001010011111110010001100011111111001011000101111000000001110010001000101011101111001111110011001100110110101001111001100001100111000110010100110000101001000010011000010111111001001110010101111010000101000011000111100000111010110011000111101100100010101000010001110111000111011101011101010111110001111010010101110100000110011001001000010111111101011110111111011010011110111100000001000000110100111100011111110000110111101000111001000010010110010011011101011100100100000;
assign EM[62] = 1024'b0001011110001111000010001001110100110110010100101011100000010000010110101000001100001111000101000000010111100011011000101100100010011101010101011000001111110111100110111111100111001100101110100011111110000000000010100110110101110011111101100001001110100010110110100000101011110101010000011010011100101001000010001111111100101110011100111000011011010111100101001001101110001110111100010110011000011000111110100000011001101101111010100000010111100010011101011001110101010011011000101100011101100101000100011101010100111001000100000000110100000111000010000010100110110101010110100110111101110110001101101010010010001001011110011000001101110110101111101101001110101000001011001011010010010111100110011011111111001100001000110110001001000111100011110111101001111110001101110011101110001001101000111101011111100111011100000111100000101101111100001111100101011111000000010001010000110111111101011011001100001011001010011010010101111100100010110001100011100001000110101000100011001110010001010110000110101001101010001111110110000111;
assign EM[63] = 1024'b0110001000101111111000001001110111010010111010101110010001001101001011111100001000001011110111010111000100100011001100100101000000111011110110101011101111010100000011110100111111110101011010111011111100110010110000101010100101000110000001011010000101010011100100100000011110110101111000010110110111110000011000101001110101110010110101101000110110010111101100111110001001100110100011001110101101110100000010010010101010001000011000001100111100010100011000000101010111111101000010011111011011101101101110100001010001100111011011110001110011101111001011010110100110100100111011010001111000001001001111000001011100101110110010010001101111010110100011000000000011011001101010011101100001110110001100110010101111110010110000010011101111110101110010101001111101100000011101111100110000000101101001001010001111001111100101100110100001101100000111110111101011110001101111100000111011100001000010000101000110101011110001001000010001111101010100100110110001110010010101100010011000010110000011000010111100010000101001000101001111011001;

genvar i;
generate
for (i=0;i<E;i=i+1) begin
    assign bind_outputs[i] = EM[i]^LBP_hvs[i];
end
endgenerate

endmodule

module BUNDLING_SPACE # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk_i,
    input  arst_n_in,
    input  [E-1:0][0:D-1] bind_outputs,
    output logic bundled_hv [0:D-1]
);

logic [E-1:0] bound_hvs [0:D-1];
logic signed [4:0] counter_array_space [0:D-1]; //maxima are 01111 and 10000

//By switching the packed and unpacked parts, can have very simple OR-tree module
genvar i10,i11;
generate
for (i11=0;i11<D/vector_fold_factor;i11=i11+1) begin
for (i10=0;i10<E/channel_fold_factor;i10=i10+1) begin
    assign bound_hvs[i11][i10] = bind_outputs[i10][i11];
end
end
endgenerate


//Bundle in space
genvar ix;
generate
for (ix=0;ix<D;ix=ix+1) begin
    adder_tree_2_directional # ( .NB_INPUTS(E) ) adder_tree_space ( .input_data(bound_hvs[ix]), .output_data(counter_array_space[ix]) );
end
endgenerate

integer iy;
always_comb begin
    for (iy=0;iy<D;iy=iy+1) begin
	bundled_hv[iy] = (counter_array_space[iy] > 0); //0 is the threshold because, this module uses the bidirectional saturating counters from the dense HDC optimizations
    end
end


endmodule


module BUNDLING_TIME # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk_i,
    input  arst_n_in,
    input  bundled_hv [0:D-1],
    output reg [0:D-1] result_hv,
    output logic [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time,
    output logic signed [4:0] counter_array [0:D-1]
);




integer i15,j2,j3,j4;
always @(posedge clk_i) begin
    for (i15=0;i15<D;i15=i15+1) begin
	if (arst_n_in == 0) begin
	    counter_bund_time <= 9'd0;
	    counter_array[i15] <= 8'd0;
	end
	else if (counter_bund_time == NB_TO_BUNDLE_IN_TIME) begin
	    counter_array[i15] <= (bundled_hv[i15]==1) ? 5'b00001:5'b11111;
	    counter_bund_time <= 1;
	end
	else if ((counter_array[i15] == 5'b01111) & (bundled_hv[i15]==1)) begin
	    counter_array[i15] <= counter_array[i15];
	    counter_bund_time <= counter_bund_time+1;
	end
	else if ((counter_array[i15] == 5'b10000) & (bundled_hv[i15]==0)) begin
	    counter_array[i15] <= counter_array[i15];
	    counter_bund_time <= counter_bund_time+1;
	end
        else begin
            counter_array[i15] <= (bundled_hv[i15]==1) ? counter_array[i15]+1:counter_array[i15]-1;
	    counter_bund_time <= counter_bund_time+1;
	end
    end
end


genvar i20;
generate
for (i20=0;i20<D;i20=i20+1) begin
always @(posedge clk_i) begin
    if (counter_bund_time == 256) begin
	result_hv[i20] <= (counter_array[i20] > 0) ? (1'b1):(1'b0); 
    end
end
end
endgenerate

endmodule


module SIMILARITY_SEARCH # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer NB_CLASSES = 2,
    parameter integer vector_fold_factor = 1, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk_i,
    input  arst_n_in,
    input  [0:D-1] result_hv,
    input  [0:D-1] ictal_hv,
    input  [0:D-1] interictal_hv,
    input  [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time,
    output classification,
    output classification_ready,
    output [$clog2(D):0] ictal_sim,
    output [$clog2(D):0] interictal_sim
);

logic [0:D-1] sim_vector;
logic [$clog2(D):0] sim_score;
logic [$clog2(D):0] sim_score_saved;
assign interictal_sim = sim_score_saved;
assign ictal_sim = sim_score;
logic [$clog2(NB_CLASSES):0] sim_counter;


always_comb begin
    if (sim_counter == 0) begin
	sim_vector = result_hv ^ interictal_hv;
    end
    else if (sim_counter == 1) begin
	sim_vector = result_hv ^ ictal_hv;
    end
end
adder_tree # ( .NB_INPUTS(D) ) adder_tree0 ( .input_data(sim_vector), .output_data(sim_score) );

always @(posedge clk_i) begin
    if (counter_bund_time == NB_TO_BUNDLE_IN_TIME) begin
	sim_counter <= 0;
    end
    else if (sim_counter == 0) begin
	sim_score_saved <= sim_score;
	sim_counter <= 1;
    end
    else if (sim_counter == 1) begin
	sim_counter <= 2;
    end
end
assign classification = (sim_score > sim_score_saved) ? 1 : 0;
assign classification_ready = (sim_counter == 1) ? 1 : 0;

endmodule


module select_if_shift # (
    parameter LENGTH_SEGMENT = 128,
    parameter SHIFT = 1
)
(
    input  [LENGTH_SEGMENT-1:0] segment,
    input  enable,
    output [LENGTH_SEGMENT-1:0] result
);
logic [LENGTH_SEGMENT-1:0] temp;
assign result = (enable) ? temp : segment;

always_comb begin
    temp[LENGTH_SEGMENT-1:SHIFT] = segment[LENGTH_SEGMENT-1-SHIFT:0];
    temp[SHIFT-1:0] = segment[LENGTH_SEGMENT-1:LENGTH_SEGMENT-SHIFT];
end

endmodule


module OR_tree # (
    parameter D = 1024,
    parameter NB_INPUTS = 64
)
(
    input [NB_INPUTS-1:0] input_hvs [D-1:0],
    output output_hv [D-1:0]
);

genvar i;
generate 
for (i=0;i<D;i=i+1) begin
    assign output_hv[i] = |input_hvs[i];
end
endgenerate 

endmodule

module adder_tree # (
    parameter NB_INPUTS,
    parameter NB_STAGES = $clog2(NB_INPUTS)
)
(
    input logic [NB_INPUTS-1:0] input_data,
    output logic [NB_STAGES:0] output_data
);

logic [NB_STAGES-1:0][(NB_INPUTS/2)-1:0][NB_STAGES:0] data; //3th part is output_data_width

genvar stage_nb, adder_nb;
generate
for (stage_nb=0;stage_nb<NB_STAGES;stage_nb=stage_nb+1) begin: stage_gen
    localparam nb_outputs_stage = NB_INPUTS >> (stage_nb+1);
    localparam data_width_stage = stage_nb+2;

    if (stage_nb == 0) begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: first_adder_gen
	    always_comb begin
		data[stage_nb][adder_nb][data_width_stage-1:0] = input_data[adder_nb*2] + input_data[adder_nb*2+1];
	    end
	end
    end
    else begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: adder_gen
	    always_comb begin
		data[stage_nb][adder_nb][data_width_stage-1:0] = 
			data[stage_nb-1][adder_nb*2][(data_width_stage-1)-1:0] + 
			data[stage_nb-1][adder_nb*2+1][(data_width_stage-1)-1:0];
	    end
        end
    end
end
endgenerate

assign output_data = data[NB_STAGES-1][0];

endmodule


module adder_tree_2_directional # (
    parameter NB_INPUTS,
    parameter NB_STAGES = $clog2(NB_INPUTS)
)
(
    input logic [NB_INPUTS-1:0] input_data,
    output logic signed [4:0] output_data
);

logic signed [NB_STAGES-1:0][(NB_INPUTS/2)-1:0][4:0] data; //3th part is output_data_width

genvar stage_nb, adder_nb;
generate
for (stage_nb=0;stage_nb<NB_STAGES;stage_nb=stage_nb+1) begin: stage_gen
    localparam nb_outputs_stage = NB_INPUTS >> (stage_nb+1);
    localparam data_width_stage = 5;

    if (stage_nb == 0) begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: first_adder_gen
	    always_comb begin
		//data[stage_nb][adder_nb][data_width_stage-1:0] = input_data[adder_nb*2] + input_data[adder_nb*2+1];
		if (input_data[adder_nb*2] == 0) begin
		    if (input_data[adder_nb*2+1] == 0) begin
			data[stage_nb][adder_nb][data_width_stage-1:0] = -2;
		    end
		    else begin
			data[stage_nb][adder_nb][data_width_stage-1:0] = 0;
		    end
		end
		else begin // == 1
		    if (input_data[adder_nb*2+1] == 0) begin
			data[stage_nb][adder_nb][data_width_stage-1:0] = 0;
		    end
		    else begin
			data[stage_nb][adder_nb][data_width_stage-1:0] = 2;
		    end
		end
	    end
	end
    end
    else begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: adder_gen
	    always_comb begin
		//data[stage_nb][adder_nb][data_width_stage-1:0] = 
			//data[stage_nb-1][adder_nb*2][(data_width_stage-1):0] + 
			//data[stage_nb-1][adder_nb*2+1][(data_width_stage-1):0];
		if (data[stage_nb-1][adder_nb*2] > 0 & data[stage_nb-1][adder_nb*2+1] > 0 & (data[stage_nb-1][adder_nb*2][(data_width_stage-1):0] + 
			data[stage_nb-1][adder_nb*2+1][(data_width_stage-1):0]) < 0) begin
		    data[stage_nb][adder_nb][data_width_stage-1:0] = 5'b01111;
		end
		else if (data[stage_nb-1][adder_nb*2] < 0 & data[stage_nb-1][adder_nb*2+1] < 0 & (data[stage_nb-1][adder_nb*2][(data_width_stage-1):0] + 
			data[stage_nb-1][adder_nb*2+1][(data_width_stage-1):0]) > 0) begin
		    data[stage_nb][adder_nb][data_width_stage-1:0] = 5'b10000;
		end
		else begin
		    data[stage_nb][adder_nb][data_width_stage-1:0] = data[stage_nb-1][adder_nb*2][(data_width_stage-1):0] + 
			data[stage_nb-1][adder_nb*2+1][(data_width_stage-1):0];
		end
	    end
        end
    end
end
endgenerate

assign output_data = data[NB_STAGES-1][0];

endmodule
