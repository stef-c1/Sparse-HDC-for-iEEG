module shift_binding_VF # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125, //0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer LBP_LENGTH = 6,
    parameter integer NB_CLASSES = 2,
    parameter integer vector_fold_factor = 2, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  [LBP_LENGTH-1:0] LBP_codes63,
    input  [LBP_LENGTH-1:0] LBP_codes62,
    input  [LBP_LENGTH-1:0] LBP_codes61,
    input  [LBP_LENGTH-1:0] LBP_codes60,
    input  [LBP_LENGTH-1:0] LBP_codes59,
    input  [LBP_LENGTH-1:0] LBP_codes58,
    input  [LBP_LENGTH-1:0] LBP_codes57,
    input  [LBP_LENGTH-1:0] LBP_codes56,
    input  [LBP_LENGTH-1:0] LBP_codes55,
    input  [LBP_LENGTH-1:0] LBP_codes54,
    input  [LBP_LENGTH-1:0] LBP_codes53,
    input  [LBP_LENGTH-1:0] LBP_codes52,
    input  [LBP_LENGTH-1:0] LBP_codes51,
    input  [LBP_LENGTH-1:0] LBP_codes50,
    input  [LBP_LENGTH-1:0] LBP_codes49,
    input  [LBP_LENGTH-1:0] LBP_codes48,
    input  [LBP_LENGTH-1:0] LBP_codes47,
    input  [LBP_LENGTH-1:0] LBP_codes46,
    input  [LBP_LENGTH-1:0] LBP_codes45,
    input  [LBP_LENGTH-1:0] LBP_codes44,
    input  [LBP_LENGTH-1:0] LBP_codes43,
    input  [LBP_LENGTH-1:0] LBP_codes42,
    input  [LBP_LENGTH-1:0] LBP_codes41,
    input  [LBP_LENGTH-1:0] LBP_codes40,
    input  [LBP_LENGTH-1:0] LBP_codes39,
    input  [LBP_LENGTH-1:0] LBP_codes38,
    input  [LBP_LENGTH-1:0] LBP_codes37,
    input  [LBP_LENGTH-1:0] LBP_codes36,
    input  [LBP_LENGTH-1:0] LBP_codes35,
    input  [LBP_LENGTH-1:0] LBP_codes34,
    input  [LBP_LENGTH-1:0] LBP_codes33,
    input  [LBP_LENGTH-1:0] LBP_codes32,
    input  [LBP_LENGTH-1:0] LBP_codes31,
    input  [LBP_LENGTH-1:0] LBP_codes30,
    input  [LBP_LENGTH-1:0] LBP_codes29,
    input  [LBP_LENGTH-1:0] LBP_codes28,
    input  [LBP_LENGTH-1:0] LBP_codes27,
    input  [LBP_LENGTH-1:0] LBP_codes26,
    input  [LBP_LENGTH-1:0] LBP_codes25,
    input  [LBP_LENGTH-1:0] LBP_codes24,
    input  [LBP_LENGTH-1:0] LBP_codes23,
    input  [LBP_LENGTH-1:0] LBP_codes22,
    input  [LBP_LENGTH-1:0] LBP_codes21,
    input  [LBP_LENGTH-1:0] LBP_codes20,
    input  [LBP_LENGTH-1:0] LBP_codes19,
    input  [LBP_LENGTH-1:0] LBP_codes18,
    input  [LBP_LENGTH-1:0] LBP_codes17,
    input  [LBP_LENGTH-1:0] LBP_codes16,
    input  [LBP_LENGTH-1:0] LBP_codes15,
    input  [LBP_LENGTH-1:0] LBP_codes14,
    input  [LBP_LENGTH-1:0] LBP_codes13,
    input  [LBP_LENGTH-1:0] LBP_codes12,
    input  [LBP_LENGTH-1:0] LBP_codes11,
    input  [LBP_LENGTH-1:0] LBP_codes10,
    input  [LBP_LENGTH-1:0] LBP_codes9,
    input  [LBP_LENGTH-1:0] LBP_codes8,
    input  [LBP_LENGTH-1:0] LBP_codes7,
    input  [LBP_LENGTH-1:0] LBP_codes6,
    input  [LBP_LENGTH-1:0] LBP_codes5,
    input  [LBP_LENGTH-1:0] LBP_codes4,
    input  [LBP_LENGTH-1:0] LBP_codes3,
    input  [LBP_LENGTH-1:0] LBP_codes2,
    input  [LBP_LENGTH-1:0] LBP_codes1,
    input  [LBP_LENGTH-1:0] LBP_codes0,
    input  [0:D-1] ictal_hv_in,
    input  [0:D-1] interictal_hv_in,
    output classification_ready,
    output [$clog2(NB_CLASSES)-1:0] classification,
    output send_next_LBP,
    output [$clog2(D):0] ictal_sim,
    output [$clog2(D):0] interictal_sim,
    output [0:D-1] result_hv2,
    output bundled_hv2 [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1],
    output [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1] bind_outputs0,
    output [(NB_SEGMENTS/vector_fold_factor)-1:0][$clog2(LENGTH_SEGMENT)-1:0] LBP_hvs0,
    output logic [$clog2(NB_TO_BUNDLE_IN_TIME)-1:0] counter_array [0:D-1],
    output logic [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time
);

//LBP_codes
logic [LBP_LENGTH-1:0] LBP_codes [E-1:0];
assign LBP_codes[63] = LBP_codes63;
assign LBP_codes[62] = LBP_codes62;
assign LBP_codes[61] = LBP_codes61;
assign LBP_codes[60] = LBP_codes60;
assign LBP_codes[59] = LBP_codes59;
assign LBP_codes[58] = LBP_codes58;
assign LBP_codes[57] = LBP_codes57;
assign LBP_codes[56] = LBP_codes56;
assign LBP_codes[55] = LBP_codes55;
assign LBP_codes[54] = LBP_codes54;
assign LBP_codes[53] = LBP_codes53;
assign LBP_codes[52] = LBP_codes52;
assign LBP_codes[51] = LBP_codes51;
assign LBP_codes[50] = LBP_codes50;
assign LBP_codes[49] = LBP_codes49;
assign LBP_codes[48] = LBP_codes48;
assign LBP_codes[47] = LBP_codes47;
assign LBP_codes[46] = LBP_codes46;
assign LBP_codes[45] = LBP_codes45;
assign LBP_codes[44] = LBP_codes44;
assign LBP_codes[43] = LBP_codes43;
assign LBP_codes[42] = LBP_codes42;
assign LBP_codes[41] = LBP_codes41;
assign LBP_codes[40] = LBP_codes40;
assign LBP_codes[39] = LBP_codes39;
assign LBP_codes[38] = LBP_codes38;
assign LBP_codes[37] = LBP_codes37;
assign LBP_codes[36] = LBP_codes36;
assign LBP_codes[35] = LBP_codes35;
assign LBP_codes[34] = LBP_codes34;
assign LBP_codes[33] = LBP_codes33;
assign LBP_codes[32] = LBP_codes32;
assign LBP_codes[31] = LBP_codes31;
assign LBP_codes[30] = LBP_codes30;
assign LBP_codes[29] = LBP_codes29;
assign LBP_codes[28] = LBP_codes28;
assign LBP_codes[27] = LBP_codes27;
assign LBP_codes[26] = LBP_codes26;
assign LBP_codes[25] = LBP_codes25;
assign LBP_codes[24] = LBP_codes24;
assign LBP_codes[23] = LBP_codes23;
assign LBP_codes[22] = LBP_codes22;
assign LBP_codes[21] = LBP_codes21;
assign LBP_codes[20] = LBP_codes20;
assign LBP_codes[19] = LBP_codes19;
assign LBP_codes[18] = LBP_codes18;
assign LBP_codes[17] = LBP_codes17;
assign LBP_codes[16] = LBP_codes16;
assign LBP_codes[15] = LBP_codes15;
assign LBP_codes[14] = LBP_codes14;
assign LBP_codes[13] = LBP_codes13;
assign LBP_codes[12] = LBP_codes12;
assign LBP_codes[11] = LBP_codes11;
assign LBP_codes[10] = LBP_codes10;
assign LBP_codes[9] = LBP_codes9;
assign LBP_codes[8] = LBP_codes8;
assign LBP_codes[7] = LBP_codes7;
assign LBP_codes[6] = LBP_codes6;
assign LBP_codes[5] = LBP_codes5;
assign LBP_codes[4] = LBP_codes4;
assign LBP_codes[3] = LBP_codes3;
assign LBP_codes[2] = LBP_codes2;
assign LBP_codes[1] = LBP_codes1;
assign LBP_codes[0] = LBP_codes0;



logic [$clog2(vector_fold_factor):0] vf_counter;

//counters for vector folding and channel folding
always @(posedge clk) begin
    if ((arst_n_in == 0) | (vector_fold_factor == 1)) begin
        vf_counter <= 'd0;
    end
    else if (vf_counter == (vector_fold_factor)) begin
        vf_counter <= 'd0;
    end
    else begin
	vf_counter <= vf_counter+1;
    end
end

//signal that need next LBP_codes
assign send_next_LBP = (vf_counter == (vector_fold_factor)) ? 1:0;


logic [LBP_LENGTH-1:0] LBP_codes_saved [E-1:0];
logic [LBP_LENGTH-1:0] LBP_codes_current [E-1:0];
//regs for LBP_values, needed if channel or vector folding is used
int i;
always_comb begin
    if (vf_counter > 0) begin
        for (i=0;i<E;i=i+1) begin
            LBP_codes_current[i] = LBP_codes_saved[i];
        end
    end
    else begin
        for (i=0;i<E;i=i+1) begin
            LBP_codes_current[i] = LBP_codes[i];
        end
    end
end

int i2;
always @(posedge clk) begin
for (i2=0;i2<E;i2=i2+1) begin
    if (arst_n_in == 0) begin
        LBP_codes_saved[i2] <= 'd0;
    end
    else begin
        LBP_codes_saved[i2] <= (vf_counter == 0) ? LBP_codes[i2]:LBP_codes_saved[i2];
    end
end
end


logic [E-1:0][$clog2(LENGTH_SEGMENT)-1:0] LBP_hvs;
//assign LBP_hvs0 = LBP_hvs[0];

logic [E-1:0][0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1] bind_outputs;
assign bind_outputs0 = bind_outputs[18];

logic bundled_hv [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1];
assign bundled_hv2 = bundled_hv;

logic [0:D-1] result_hv;
//assign result_hv2 = result_hv;
//logic [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time;
//logic [$clog2(NB_TO_BUNDLE_IN_TIME)-1:0] counter_array [0:D-1];

logic [0:D-1] ictal_hv;
logic [0:D-1] interictal_hv;


assign ictal_hv = (arst_n_in) ? ictal_hv : ictal_hv_in;
assign interictal_hv = (arst_n_in) ? interictal_hv : interictal_hv_in;

//The Big Five
IM #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
IM_module (.clk(clk), .arst_n_in(arst_n_in), .LBP_codes(LBP_codes_current), .vf_counter(vf_counter), .LBP_hvs(LBP_hvs));

BINDING2 #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BINDING_module (.clk(clk), .arst_n_in(arst_n_in), .LBP_hvs(LBP_hvs), .vf_counter(vf_counter), .bind_outputs(bind_outputs));

BUNDLING_SPACE2 #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BUNDLING_SPACE_module (.clk(clk), .arst_n_in(arst_n_in), .bind_outputs(bind_outputs), .vf_counter(vf_counter), .bundled_hv_e(bundled_hv));

BUNDLING_TIME #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .NB_TO_BUNDLE_IN_TIME(NB_TO_BUNDLE_IN_TIME), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor)) 
BUNDLING_TIME_module (.clk(clk), .arst_n_in(arst_n_in), .bundled_hv(bundled_hv), .vf_counter(vf_counter), .result_hv(result_hv), .counter_bund_time(counter_bund_time), .counter_array(counter_array));

SIMILARITY_SEARCH #(.D(D), /*.p_sparse(p_sparse),*/ .E(E), .NB_SEGMENTS(NB_SEGMENTS), .LENGTH_SEGMENT(LENGTH_SEGMENT), .NB_TO_BUNDLE_IN_TIME(NB_TO_BUNDLE_IN_TIME), .LBP_LENGTH(LBP_LENGTH), .vector_fold_factor(vector_fold_factor), .channel_fold_factor(channel_fold_factor), .NB_CLASSES(NB_CLASSES)) 
SIMILARITY_SEARCH_module (.clk(clk), .arst_n_in(arst_n_in), .result_hv(result_hv), .ictal_hv(ictal_hv), .interictal_hv(interictal_hv), .vf_counter(vf_counter), .counter_bund_time(counter_bund_time), .classification(classification), .classification_ready(classification_ready), .ictal_sim(ictal_sim), .interictal_sim(interictal_sim));


endmodule


module IM # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 4, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  [LBP_LENGTH-1:0] LBP_codes [E-1:0],
    input  [$clog2(vector_fold_factor):0] vf_counter,
    output logic [E/channel_fold_factor-1:0][$clog2(LENGTH_SEGMENT)-1:0] LBP_hvs
);

genvar i,j;
generate
for (i=0;i<E;i=i+1) begin
    assign LBP_hvs[i] = {1'b0,LBP_codes[i]};
end
endgenerate

endmodule

module BINDING2 # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 4, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  [E-1:0][$clog2(LENGTH_SEGMENT)-1:0] LBP_hvs,
    input  [$clog2(vector_fold_factor):0] vf_counter,
    output [E-1:0][0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1] bind_outputs

);
logic [$clog2(LENGTH_SEGMENT):0][E-1:0][0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1] intermediate_bind_outputs;
assign bind_outputs = intermediate_bind_outputs[$clog2(LENGTH_SEGMENT)-1];


logic [E-1:0][0:LENGTH_SEGMENT*NB_SEGMENTS-1] EM;

assign EM[0] = 1024'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
assign EM[1] = 1024'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
assign EM[2] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
assign EM[3] = 1024'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[4] = 1024'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[5] = 1024'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
assign EM[6] = 1024'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
assign EM[7] = 1024'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
assign EM[8] = 1024'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
assign EM[9] = 1024'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
assign EM[10] = 1024'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[11] = 1024'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[12] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
assign EM[13] = 1024'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[14] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
assign EM[15] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
assign EM[16] = 1024'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
assign EM[17] = 1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[18] = 1024'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[19] = 1024'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
assign EM[20] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
assign EM[21] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[22] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
assign EM[23] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[24] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
assign EM[25] = 1024'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[26] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[27] = 1024'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
assign EM[28] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[29] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[30] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
assign EM[31] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
assign EM[32] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[33] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
assign EM[34] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[35] = 1024'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[36] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[37] = 1024'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
assign EM[38] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
assign EM[39] = 1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
assign EM[40] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[41] = 1024'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
assign EM[42] = 1024'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
assign EM[43] = 1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[44] = 1024'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[45] = 1024'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[46] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
assign EM[47] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
assign EM[48] = 1024'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
assign EM[49] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
assign EM[50] = 1024'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
assign EM[51] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
assign EM[52] = 1024'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[53] = 1024'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[54] = 1024'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[55] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[56] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
assign EM[57] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[58] = 1024'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[59] = 1024'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
assign EM[60] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
assign EM[61] = 1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
assign EM[62] = 1024'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign EM[63] = 1024'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

//set EM as inputs to the binding
integer k,k50,k_cf;
always_comb begin
for (k=0;k<vector_fold_factor;k=k+1) begin
for (k50=0;k50<E;k50=k50+1) begin
    if (vf_counter === 0) begin //if (vf_counter == 0)
        intermediate_bind_outputs[0][k50] = EM[k50][(vector_fold_factor-1)*NB_SEGMENTS/vector_fold_factor*LENGTH_SEGMENT +: NB_SEGMENTS/vector_fold_factor*LENGTH_SEGMENT];
    end
    else if (vf_counter === k+1) begin
        intermediate_bind_outputs[0][k50] = EM[k50][k*NB_SEGMENTS/vector_fold_factor*LENGTH_SEGMENT +: NB_SEGMENTS/vector_fold_factor*LENGTH_SEGMENT];
    end
end
end
end


reg [E-1:0][2**(LBP_LENGTH)-1:0] to_slide_in_reg; 
wire [E-1:0][2**(LBP_LENGTH)-1:0] to_slide_in_reg_input; 

always @(posedge clk) begin
    if (arst_n_in == 0)
	to_slide_in_reg <= 'd0;
    else
	to_slide_in_reg <= to_slide_in_reg_input;
end


//All the E/channel_fold_factor*NB_SEGMENTS/vector_fold_factor binding units
genvar i2,i4;
generate 
  if (vector_fold_factor == 1) begin
    for (i4=0;i4<E/channel_fold_factor;i4=i4+1) begin: binding_i4_gen
    for (i2=0;i2<LBP_LENGTH;i2=i2+1) begin: binding_i2_gen
	select_if_shift #(.LENGTH_SEGMENT(LENGTH_SEGMENT*NB_SEGMENTS),.SHIFT(2**(i2))) select_if_shift0 (.segment(intermediate_bind_outputs[i2][i4]), .enable(LBP_hvs[i4][i2]), .result(intermediate_bind_outputs[i2+1][i4]));
    end
    end
  end
  else begin
    for (i4=0;i4<E/channel_fold_factor;i4=i4+1) begin: binding_i4_gen
    for (i2=0;i2<LBP_LENGTH;i2=i2+1) begin: binding_i2_gen
	select_if_shift2 #(.LENGTH_SEGMENT(LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor),.SHIFT(2**(i2))) select_if_shift02 (.segment(intermediate_bind_outputs[i2][i4]), .enable(LBP_hvs[i4][i2]), .to_slide_in(to_slide_in_reg[i4][(2**(i2)-1) +: 2**(i2)]), .result(intermediate_bind_outputs[i2+1][i4]), .to_slide_out(to_slide_in_reg_input[i4][(2**(i2)-1) +: 2**(i2)]));
    end
    end
  end
endgenerate

endmodule

module BUNDLING_SPACE2 # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 4, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  [E-1:0][0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1] bind_outputs,
    input  [$clog2(vector_fold_factor):0] vf_counter,
    output bundled_hv_e [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1]
);

logic [E-1:0] bound_hvs [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1];
logic bundled_hv_e2 [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1];


genvar i88;
generate
for (i88=0;i88<D/vector_fold_factor;i88=i88+1) begin
assign bundled_hv_e[i88] = (vf_counter === 0) ? 'd0:bundled_hv_e2[i88];
end
endgenerate

//By switching the packed and unpacked parts, can have very simple OR-tree module
genvar i10,i11;
generate
for (i11=0;i11<D/vector_fold_factor;i11=i11+1) begin
for (i10=0;i10<E;i10=i10+1) begin
    assign bound_hvs[i11][i10] = bind_outputs[i10][i11];
end
end
endgenerate


//Bundle in space
OR_tree #(.D(D/vector_fold_factor),.NB_INPUTS(E)) OR_tree0 (.input_hvs(bound_hvs), .output_hv(bundled_hv_e2));


endmodule


module BUNDLING_TIME # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer vector_fold_factor = 4, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  bundled_hv [0:LENGTH_SEGMENT*NB_SEGMENTS/vector_fold_factor-1],
    input  [$clog2(vector_fold_factor):0] vf_counter,
    output logic [0:D-1] result_hv,
    output logic [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time,
    output logic [$clog2(NB_TO_BUNDLE_IN_TIME)-1:0] counter_array [0:D-1]
);

//logic [$clog2(NB_TO_BUNDLE_IN_TIME)-1:0] counter_array [0:D-1];



integer i15,j2,j3,j4;
always @(posedge clk) begin
    for (i15=0;i15<D/vector_fold_factor;i15=i15+1) begin
	if (arst_n_in == 0) begin
	    counter_bund_time <= 9'd0;//'0
	    counter_array[i15] <= 8'd0;//'0;
            for (j4=1;j4<vector_fold_factor;j4=j4+1) begin
		counter_array[i15+j4*D/vector_fold_factor] <= 8'd0;//'0;
	    end
	end
	else if (counter_bund_time == NB_TO_BUNDLE_IN_TIME) begin
            for (j3=0;j3<vector_fold_factor;j3=j3+1) begin
		if (vf_counter === (j3+1)) begin
		    counter_array[i15+j3*D/vector_fold_factor] <= bundled_hv[i15];
		    if (vf_counter === (vector_fold_factor)) begin
			counter_bund_time <= 1;
		    end
		end
	    end
	end
	else begin
    	    for (j2=0;j2<vector_fold_factor;j2=j2+1) begin
	        if (vf_counter === (j2+1)) begin
                    counter_array[i15+j2*D/vector_fold_factor] <= (bundled_hv[i15]===1) ? counter_array[i15+j2*D/vector_fold_factor]+1:counter_array[i15+j2*D/vector_fold_factor];
	        end
	    end
	    counter_bund_time <= (vf_counter === (vector_fold_factor)) ? counter_bund_time+1:counter_bund_time;
	end
    end
end


genvar i20;
generate
for (i20=0;i20<D;i20=i20+1) begin
always @(posedge clk) begin
    if ((counter_bund_time == NB_TO_BUNDLE_IN_TIME) & (vf_counter === 0)) begin
	result_hv[i20] <= (counter_array[i20] > 8'h82) ? (1'b1):(1'b0); //h82
    end
end
end
endgenerate

endmodule


module SIMILARITY_SEARCH # (
    parameter integer D = 1024,
    //parameter real p_sparse = 0.0078125,
    parameter integer E = 64,
    parameter integer NB_TO_BUNDLE_IN_TIME = 256,
    parameter integer NB_SEGMENTS = 8,
    parameter integer LENGTH_SEGMENT = 128,
    parameter integer LBP_LENGTH = 6,
    parameter integer NB_CLASSES = 2,
    parameter integer vector_fold_factor = 4, //either 1,2,4...NB_SEGMENTS
    parameter integer channel_fold_factor = 1 //either 1,2,4...E (if E is a power of 2)
)
(
    input  clk,
    input  arst_n_in,
    input  [0:D-1] result_hv,
    input  [0:D-1] ictal_hv,
    input  [0:D-1] interictal_hv,
    input  [$clog2(vector_fold_factor):0] vf_counter,
    input  [$clog2(NB_TO_BUNDLE_IN_TIME):0] counter_bund_time,
    output classification,
    output classification_ready,
    output [$clog2(D):0] ictal_sim,
    output [$clog2(D):0] interictal_sim
);

logic [0:D-1] sim_vector;
logic [$clog2(D):0] sim_score;
logic [$clog2(D):0] sim_score_saved;
assign interictal_sim = sim_score_saved;
assign ictal_sim = sim_score;
logic [$clog2(NB_CLASSES):0] sim_counter;


always_comb begin
    if (sim_counter == 0) begin
	sim_vector = result_hv & interictal_hv;
    end
    else if (sim_counter == 1) begin
	sim_vector = result_hv & ictal_hv;
    end
end
adder_tree # ( .NB_INPUTS(D) ) adder_tree0 ( .input_data(sim_vector), .output_data(sim_score) );

always @(posedge clk) begin
    if ((counter_bund_time == NB_TO_BUNDLE_IN_TIME) & (vf_counter == 0)) begin
	sim_counter <= 0;
    end
    else if (sim_counter == 0) begin
	sim_score_saved <= sim_score;
	sim_counter <= 1;
    end
    else if (sim_counter == 1) begin
	sim_counter <= 2;
    end
end
assign classification = (sim_score > sim_score_saved) ? 1 : 0;
assign classification_ready = (sim_counter == 1) ? 1 : 0;

endmodule


module select_if_shift # (
    parameter LENGTH_SEGMENT = 128,
    parameter SHIFT = 1
)
(
    input  [LENGTH_SEGMENT-1:0] segment,
    input  enable,
    output [LENGTH_SEGMENT-1:0] result
);
logic [LENGTH_SEGMENT-1:0] temp;
assign result = (enable) ? temp : segment;

always_comb begin
    temp[LENGTH_SEGMENT-1:SHIFT] = segment[LENGTH_SEGMENT-1-SHIFT:0];
    temp[SHIFT-1:0] = segment[LENGTH_SEGMENT-1:LENGTH_SEGMENT-SHIFT];
end

endmodule

module select_if_shift2 # (
    parameter LENGTH_SEGMENT = 1024,
    parameter SHIFT = 1
)
(
    input  [0:LENGTH_SEGMENT-1] segment,
    input  [0:SHIFT-1] to_slide_in,
    input  enable,
    output [0:LENGTH_SEGMENT-1] result,
    output logic [0:SHIFT-1] to_slide_out
);
logic [0:LENGTH_SEGMENT-1] temp;
assign result = (enable) ? temp : segment;

always_comb begin
    temp[SHIFT:LENGTH_SEGMENT-1] = segment[0:LENGTH_SEGMENT-1-SHIFT];
    temp[0:SHIFT-1] = to_slide_in;
    to_slide_out = segment[LENGTH_SEGMENT-SHIFT:LENGTH_SEGMENT-1];
end

endmodule

/*module select_if_shift2 # ( //Needs to shift oppositely!!!
    parameter LENGTH_SEGMENT = 1024,
    parameter SHIFT = 1
)
(
    input  [LENGTH_SEGMENT-1:0] segment,
    input  [SHIFT-1:0] to_slide_in,
    input  enable,
    output [LENGTH_SEGMENT-1:0] result,
    output logic [SHIFT-1:0] to_slide_out
);
logic [LENGTH_SEGMENT-1:0] temp;
assign result = (enable) ? temp : segment;

always_comb begin
    temp[LENGTH_SEGMENT-1:SHIFT] = segment[LENGTH_SEGMENT-1-SHIFT:0];
    temp[SHIFT-1:0] = to_slide_in;
    to_slide_out = segment[LENGTH_SEGMENT-1:LENGTH_SEGMENT-SHIFT];
end

endmodule
*/

module OR_tree # (
    parameter D = 1024,
    parameter NB_INPUTS = 64
)
(
    input [NB_INPUTS-1:0] input_hvs [D-1:0],
    output output_hv [D-1:0]
);

genvar i;
generate 
for (i=0;i<D;i=i+1) begin
    assign output_hv[i] = |input_hvs[i];
end
endgenerate 

endmodule

module adder_tree # (
    parameter NB_INPUTS,
    parameter NB_STAGES = $clog2(NB_INPUTS)
)
(
    input logic [NB_INPUTS-1:0] input_data,
    output logic [NB_STAGES:0] output_data
);

logic [NB_STAGES-1:0][(NB_INPUTS/2)-1:0][NB_STAGES:0] data; //3th part is output_data_width

genvar stage_nb, adder_nb;
generate
for (stage_nb=0;stage_nb<NB_STAGES;stage_nb=stage_nb+1) begin: stage_gen
    localparam nb_outputs_stage = NB_INPUTS >> (stage_nb+1);
    localparam data_width_stage = stage_nb+2;

    if (stage_nb == 0) begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: first_adder_gen
	    always_comb begin
		data[stage_nb][adder_nb][data_width_stage-1:0] = input_data[adder_nb*2] + input_data[adder_nb*2+1];
	    end
	end
    end
    else begin
	for (adder_nb=0;adder_nb<nb_outputs_stage;adder_nb=adder_nb+1) begin: adder_gen
	    always_comb begin
		data[stage_nb][adder_nb][data_width_stage-1:0] = 
			data[stage_nb-1][adder_nb*2][(data_width_stage-1)-1:0] + 
			data[stage_nb-1][adder_nb*2+1][(data_width_stage-1)-1:0];
	    end
        end
    end
end
endgenerate

assign output_data = data[NB_STAGES-1][0];

endmodule
